module MCacheCtrl(
  input         clock,
  input         reset,
  output        io_fetchEna,
  output        io_ctrlrepl_wEna,
  output [31:0] io_ctrlrepl_wData,
  output [31:0] io_ctrlrepl_wAddr,
  output        io_ctrlrepl_wTag,
  output [10:0] io_ctrlrepl_addrEven,
  output [10:0] io_ctrlrepl_addrOdd,
  output        io_ctrlrepl_instrStall,
  input         io_replctrl_hit,
  input  [31:0] io_femcache_addrEven,
  input  [31:0] io_femcache_addrOdd,
  input         io_exmcache_doCallRet,
  input  [31:0] io_exmcache_callRetBase,
  output [2:0]  io_ocp_port_M_Cmd,
  output [31:0] io_ocp_port_M_Addr,
  input  [1:0]  io_ocp_port_S_Resp,
  input  [31:0] io_ocp_port_S_Data,
  input         io_ocp_port_S_CmdAccept,
  output        io_illMem,
  output        io_forceHit
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] stateReg; // @[MCache.scala 293:21]
  reg [2:0] ocpCmdReg; // @[MCache.scala 302:22]
  reg [31:0] ocpAddrReg; // @[MCache.scala 303:23]
  reg [10:0] transferSizeReg; // @[MCache.scala 305:28]
  reg [10:0] fetchCntReg; // @[MCache.scala 306:24]
  reg [1:0] burstCntReg; // @[MCache.scala 307:24]
  reg [31:0] callRetBaseReg; // @[MCache.scala 309:27]
  wire [31:0] msizeAddr = callRetBaseReg - 32'h1; // @[MCache.scala 311:34]
  reg [31:0] addrEvenReg; // @[MCache.scala 312:24]
  reg [31:0] addrOddReg; // @[MCache.scala 313:23]
  reg [1:0] ocpSlaveReg_Resp; // @[MCache.scala 315:24]
  reg [31:0] ocpSlaveReg_Data; // @[MCache.scala 315:24]
  wire [2:0] _GEN_0 = io_ocp_port_S_CmdAccept ? 3'h0 : ocpCmdReg; // @[MCache.scala 330:46 MCache.scala 331:15 MCache.scala 302:22]
  wire [33:0] _T_2 = {ocpAddrReg,2'h0}; // @[Cat.scala 30:58]
  wire  _T_5 = ~io_ocp_port_S_CmdAccept; // @[MCache.scala 359:37]
  wire [2:0] _GEN_4 = ~io_ocp_port_S_CmdAccept ? 3'h2 : _GEN_0; // @[MCache.scala 359:50 MCache.scala 360:19]
  wire [29:0] hi = msizeAddr[31:2]; // @[MCache.scala 362:42]
  wire [33:0] _T_6 = {hi,4'h0}; // @[Cat.scala 30:58]
  wire [31:0] _hi_T = {hi,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_5 = io_replctrl_hit ? io_femcache_addrEven : addrEvenReg; // @[MCache.scala 349:39 MCache.scala 350:16 MCache.scala 318:12]
  wire [31:0] _GEN_6 = io_replctrl_hit ? io_femcache_addrOdd : addrOddReg; // @[MCache.scala 349:39 MCache.scala 351:15 MCache.scala 319:11]
  wire [1:0] _GEN_7 = io_replctrl_hit ? burstCntReg : 2'h0; // @[MCache.scala 349:39 MCache.scala 307:24 MCache.scala 355:19]
  wire [2:0] _GEN_8 = io_replctrl_hit ? ocpCmdReg : 3'h2; // @[MCache.scala 349:39 MCache.scala 336:21 MCache.scala 358:25]
  wire [2:0] _GEN_9 = io_replctrl_hit ? _GEN_0 : _GEN_4; // @[MCache.scala 349:39]
  wire [33:0] _GEN_10 = io_replctrl_hit ? _T_2 : _T_6; // @[MCache.scala 349:39 MCache.scala 335:22 MCache.scala 362:26]
  wire [31:0] _GEN_11 = io_replctrl_hit ? ocpAddrReg : _hi_T; // @[MCache.scala 349:39 MCache.scala 303:23 MCache.scala 364:18]
  wire [2:0] _GEN_12 = io_replctrl_hit ? stateReg : 3'h1; // @[MCache.scala 349:39 MCache.scala 293:21 MCache.scala 367:16]
  wire [31:0] _GEN_13 = stateReg == 3'h0 ? _GEN_5 : addrEvenReg; // @[MCache.scala 348:33 MCache.scala 318:12]
  wire [31:0] _GEN_14 = stateReg == 3'h0 ? _GEN_6 : addrOddReg; // @[MCache.scala 348:33 MCache.scala 319:11]
  wire [1:0] _GEN_15 = stateReg == 3'h0 ? _GEN_7 : burstCntReg; // @[MCache.scala 348:33 MCache.scala 307:24]
  wire [2:0] _GEN_16 = stateReg == 3'h0 ? _GEN_8 : ocpCmdReg; // @[MCache.scala 348:33 MCache.scala 336:21]
  wire [2:0] _GEN_17 = stateReg == 3'h0 ? _GEN_9 : _GEN_0; // @[MCache.scala 348:33]
  wire [33:0] _GEN_18 = stateReg == 3'h0 ? _GEN_10 : _T_2; // @[MCache.scala 348:33 MCache.scala 335:22]
  wire [31:0] _GEN_19 = stateReg == 3'h0 ? _GEN_11 : ocpAddrReg; // @[MCache.scala 348:33 MCache.scala 303:23]
  wire [2:0] _GEN_20 = stateReg == 3'h0 ? _GEN_12 : stateReg; // @[MCache.scala 348:33 MCache.scala 293:21]
  wire  _T_8 = ocpSlaveReg_Resp == 2'h1; // @[MCache.scala 373:28]
  wire [1:0] _T_10 = burstCntReg + 2'h1; // @[MCache.scala 374:34]
  wire  _T_12 = burstCntReg == msizeAddr[1:0]; // @[MCache.scala 375:25]
  wire [11:0] _T_15 = ocpSlaveReg_Data[13:2] - 12'h1; // @[MCache.scala 378:33]
  wire  _T_16 = burstCntReg == 2'h3; // @[MCache.scala 380:27]
  wire [2:0] _GEN_21 = _T_5 ? 3'h2 : _GEN_17; // @[MCache.scala 382:54 MCache.scala 383:23]
  wire [33:0] _T_18 = {callRetBaseReg,2'h0}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_22 = burstCntReg == 2'h3 ? 3'h2 : _GEN_16; // @[MCache.scala 380:55 MCache.scala 381:29]
  wire [2:0] _GEN_23 = burstCntReg == 2'h3 ? _GEN_21 : _GEN_17; // @[MCache.scala 380:55]
  wire [33:0] _GEN_24 = burstCntReg == 2'h3 ? _T_18 : _GEN_18; // @[MCache.scala 380:55 MCache.scala 385:30]
  wire [31:0] _GEN_25 = burstCntReg == 2'h3 ? callRetBaseReg : _GEN_19; // @[MCache.scala 380:55 MCache.scala 386:22]
  wire [1:0] _GEN_26 = burstCntReg == 2'h3 ? 2'h0 : _T_10; // @[MCache.scala 380:55 MCache.scala 387:23 MCache.scala 374:19]
  wire [11:0] _GEN_139 = {{11'd0}, ocpSlaveReg_Data[2]}; // @[MCache.scala 392:22]
  wire [11:0] _T_21 = ocpSlaveReg_Data[13:2] + _GEN_139; // @[MCache.scala 392:22]
  wire [11:0] _GEN_27 = burstCntReg == msizeAddr[1:0] ? _T_15 : {{1'd0}, transferSizeReg}; // @[MCache.scala 375:66 MCache.scala 378:25 MCache.scala 305:28]
  wire [10:0] _GEN_28 = burstCntReg == msizeAddr[1:0] ? 11'h0 : fetchCntReg; // @[MCache.scala 375:66 MCache.scala 379:21 MCache.scala 306:24]
  wire [2:0] _GEN_29 = burstCntReg == msizeAddr[1:0] ? _GEN_22 : _GEN_16; // @[MCache.scala 375:66]
  wire [2:0] _GEN_30 = burstCntReg == msizeAddr[1:0] ? _GEN_23 : _GEN_17; // @[MCache.scala 375:66]
  wire [33:0] _GEN_31 = burstCntReg == msizeAddr[1:0] ? _GEN_24 : _GEN_18; // @[MCache.scala 375:66]
  wire [31:0] _GEN_32 = burstCntReg == msizeAddr[1:0] ? _GEN_25 : _GEN_19; // @[MCache.scala 375:66]
  wire [1:0] _GEN_33 = burstCntReg == msizeAddr[1:0] ? _GEN_26 : _T_10; // @[MCache.scala 375:66 MCache.scala 374:19]
  wire [11:0] _GEN_35 = burstCntReg == msizeAddr[1:0] ? _T_21 : 12'h0; // @[MCache.scala 375:66 MCache.scala 392:15 MCache.scala 320:9]
  wire [31:0] _GEN_36 = burstCntReg == msizeAddr[1:0] ? callRetBaseReg : 32'h0; // @[MCache.scala 375:66 MCache.scala 394:15 MCache.scala 323:9]
  wire [2:0] _GEN_37 = burstCntReg == msizeAddr[1:0] ? 3'h2 : _GEN_20; // @[MCache.scala 375:66 MCache.scala 395:18]
  wire [1:0] _GEN_38 = ocpSlaveReg_Resp == 2'h1 ? _GEN_33 : _GEN_15; // @[MCache.scala 373:45]
  wire [11:0] _GEN_39 = ocpSlaveReg_Resp == 2'h1 ? _GEN_27 : {{1'd0}, transferSizeReg}; // @[MCache.scala 373:45 MCache.scala 305:28]
  wire [10:0] _GEN_40 = ocpSlaveReg_Resp == 2'h1 ? _GEN_28 : fetchCntReg; // @[MCache.scala 373:45 MCache.scala 306:24]
  wire [2:0] _GEN_41 = ocpSlaveReg_Resp == 2'h1 ? _GEN_29 : _GEN_16; // @[MCache.scala 373:45]
  wire [2:0] _GEN_42 = ocpSlaveReg_Resp == 2'h1 ? _GEN_30 : _GEN_17; // @[MCache.scala 373:45]
  wire [33:0] _GEN_43 = ocpSlaveReg_Resp == 2'h1 ? _GEN_31 : _GEN_18; // @[MCache.scala 373:45]
  wire [31:0] _GEN_44 = ocpSlaveReg_Resp == 2'h1 ? _GEN_32 : _GEN_19; // @[MCache.scala 373:45]
  wire  _GEN_45 = ocpSlaveReg_Resp == 2'h1 & _T_12; // @[MCache.scala 373:45 MCache.scala 321:8]
  wire [11:0] _GEN_46 = ocpSlaveReg_Resp == 2'h1 ? _GEN_35 : 12'h0; // @[MCache.scala 373:45 MCache.scala 320:9]
  wire [31:0] _GEN_47 = ocpSlaveReg_Resp == 2'h1 ? _GEN_36 : 32'h0; // @[MCache.scala 373:45 MCache.scala 323:9]
  wire [2:0] _GEN_48 = ocpSlaveReg_Resp == 2'h1 ? _GEN_37 : _GEN_20; // @[MCache.scala 373:45]
  wire  _GEN_49 = stateReg == 3'h1 ? 1'h0 : 1'h1; // @[MCache.scala 371:33 MCache.scala 372:14 MCache.scala 324:12]
  wire [1:0] _GEN_50 = stateReg == 3'h1 ? _GEN_38 : _GEN_15; // @[MCache.scala 371:33]
  wire [11:0] _GEN_51 = stateReg == 3'h1 ? _GEN_39 : {{1'd0}, transferSizeReg}; // @[MCache.scala 371:33 MCache.scala 305:28]
  wire [10:0] _GEN_52 = stateReg == 3'h1 ? _GEN_40 : fetchCntReg; // @[MCache.scala 371:33 MCache.scala 306:24]
  wire [2:0] _GEN_53 = stateReg == 3'h1 ? _GEN_41 : _GEN_16; // @[MCache.scala 371:33]
  wire [2:0] _GEN_54 = stateReg == 3'h1 ? _GEN_42 : _GEN_17; // @[MCache.scala 371:33]
  wire [33:0] _GEN_55 = stateReg == 3'h1 ? _GEN_43 : _GEN_18; // @[MCache.scala 371:33]
  wire [31:0] _GEN_56 = stateReg == 3'h1 ? _GEN_44 : _GEN_19; // @[MCache.scala 371:33]
  wire [11:0] _GEN_58 = stateReg == 3'h1 ? _GEN_46 : 12'h0; // @[MCache.scala 371:33 MCache.scala 320:9]
  wire [31:0] _GEN_59 = stateReg == 3'h1 ? _GEN_47 : 32'h0; // @[MCache.scala 371:33 MCache.scala 323:9]
  wire [2:0] _GEN_60 = stateReg == 3'h1 ? _GEN_48 : _GEN_20; // @[MCache.scala 371:33]
  wire [10:0] _T_26 = fetchCntReg + 11'h1; // @[MCache.scala 405:36]
  wire [2:0] _GEN_61 = _T_5 ? 3'h2 : _GEN_54; // @[MCache.scala 411:56 MCache.scala 412:25]
  wire [31:0] _GEN_140 = {{21'd0}, fetchCntReg}; // @[MCache.scala 414:54]
  wire [31:0] _T_33 = callRetBaseReg + _GEN_140; // @[MCache.scala 414:54]
  wire [31:0] hi_1 = _T_33 + 32'h1; // @[MCache.scala 414:68]
  wire [33:0] _T_35 = {hi_1,2'h0}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_62 = _T_16 ? 3'h2 : _GEN_53; // @[MCache.scala 409:57 MCache.scala 410:31]
  wire [2:0] _GEN_63 = _T_16 ? _GEN_61 : _GEN_54; // @[MCache.scala 409:57]
  wire [33:0] _GEN_64 = _T_16 ? _T_35 : _GEN_55; // @[MCache.scala 409:57 MCache.scala 414:32]
  wire [31:0] _GEN_65 = _T_16 ? hi_1 : _GEN_56; // @[MCache.scala 409:57 MCache.scala 415:24]
  wire [31:0] _GEN_68 = _T_16 ? io_femcache_addrEven : _GEN_13; // @[MCache.scala 421:57 MCache.scala 423:22]
  wire [31:0] _GEN_69 = _T_16 ? io_femcache_addrOdd : _GEN_14; // @[MCache.scala 421:57 MCache.scala 424:21]
  wire [2:0] _GEN_70 = _T_16 ? 3'h0 : _GEN_60; // @[MCache.scala 421:57 MCache.scala 425:22]
  wire [2:0] _GEN_71 = fetchCntReg < transferSizeReg ? _GEN_62 : _GEN_53; // @[MCache.scala 407:45]
  wire [2:0] _GEN_72 = fetchCntReg < transferSizeReg ? _GEN_63 : _GEN_54; // @[MCache.scala 407:45]
  wire [33:0] _GEN_73 = fetchCntReg < transferSizeReg ? _GEN_64 : _GEN_55; // @[MCache.scala 407:45]
  wire [1:0] _GEN_75 = fetchCntReg < transferSizeReg ? _GEN_26 : _T_10; // @[MCache.scala 407:45 MCache.scala 406:21]
  wire  _GEN_76 = fetchCntReg < transferSizeReg ? 1'h0 : _T_16; // @[MCache.scala 407:45 MCache.scala 402:14]
  wire [31:0] _GEN_77 = fetchCntReg < transferSizeReg ? _GEN_13 : _GEN_68; // @[MCache.scala 407:45]
  wire [31:0] _GEN_78 = fetchCntReg < transferSizeReg ? _GEN_14 : _GEN_69; // @[MCache.scala 407:45]
  wire [2:0] _GEN_79 = fetchCntReg < transferSizeReg ? _GEN_60 : _GEN_70; // @[MCache.scala 407:45]
  wire [1:0] _GEN_81 = _T_8 ? _GEN_75 : _GEN_50; // @[MCache.scala 404:47]
  wire [2:0] _GEN_82 = _T_8 ? _GEN_71 : _GEN_53; // @[MCache.scala 404:47]
  wire [2:0] _GEN_83 = _T_8 ? _GEN_72 : _GEN_54; // @[MCache.scala 404:47]
  wire [33:0] _GEN_84 = _T_8 ? _GEN_73 : _GEN_55; // @[MCache.scala 404:47]
  wire  _GEN_86 = _T_8 & _GEN_76; // @[MCache.scala 404:47 MCache.scala 402:14]
  wire [31:0] _GEN_87 = _T_8 ? _GEN_77 : _GEN_13; // @[MCache.scala 404:47]
  wire [31:0] _GEN_88 = _T_8 ? _GEN_78 : _GEN_14; // @[MCache.scala 404:47]
  wire [2:0] _GEN_89 = _T_8 ? _GEN_79 : _GEN_60; // @[MCache.scala 404:47]
  wire [31:0] _GEN_90 = _T_8 ? ocpSlaveReg_Data : {{20'd0}, _GEN_58}; // @[MCache.scala 404:47 MCache.scala 429:15]
  wire [1:0] _GEN_92 = _T_8 ? _T_10 : _GEN_50; // @[MCache.scala 436:47 MCache.scala 437:21]
  wire [1:0] _GEN_98 = fetchCntReg <= transferSizeReg ? _GEN_81 : _GEN_92; // @[MCache.scala 403:43]
  wire [2:0] _GEN_99 = fetchCntReg <= transferSizeReg ? _GEN_82 : _GEN_53; // @[MCache.scala 403:43]
  wire [33:0] _GEN_101 = fetchCntReg <= transferSizeReg ? _GEN_84 : _GEN_55; // @[MCache.scala 403:43]
  wire  _GEN_103 = fetchCntReg <= transferSizeReg ? _GEN_86 : _T_16; // @[MCache.scala 403:43]
  wire [31:0] _GEN_104 = fetchCntReg <= transferSizeReg ? _GEN_87 : _GEN_68; // @[MCache.scala 403:43]
  wire [31:0] _GEN_105 = fetchCntReg <= transferSizeReg ? _GEN_88 : _GEN_69; // @[MCache.scala 403:43]
  wire [2:0] _GEN_106 = fetchCntReg <= transferSizeReg ? _GEN_89 : _GEN_70; // @[MCache.scala 403:43]
  wire [31:0] _GEN_107 = fetchCntReg <= transferSizeReg ? _GEN_90 : {{20'd0}, _GEN_58}; // @[MCache.scala 403:43]
  wire  _GEN_108 = fetchCntReg <= transferSizeReg & _T_8; // @[MCache.scala 403:43 MCache.scala 322:8]
  wire [31:0] _GEN_109 = fetchCntReg <= transferSizeReg ? {{21'd0}, fetchCntReg} : _GEN_59; // @[MCache.scala 403:43 MCache.scala 432:13]
  wire [1:0] _GEN_112 = stateReg == 3'h2 ? _GEN_98 : _GEN_50; // @[MCache.scala 401:37]
  wire [2:0] _GEN_113 = stateReg == 3'h2 ? _GEN_99 : _GEN_53; // @[MCache.scala 401:37]
  wire [33:0] _GEN_115 = stateReg == 3'h2 ? _GEN_101 : _GEN_55; // @[MCache.scala 401:37]
  wire [31:0] addrEven = stateReg == 3'h2 ? _GEN_104 : _GEN_13; // @[MCache.scala 401:37]
  wire [31:0] addrOdd = stateReg == 3'h2 ? _GEN_105 : _GEN_14; // @[MCache.scala 401:37]
  wire [2:0] _GEN_119 = stateReg == 3'h2 ? _GEN_106 : _GEN_60; // @[MCache.scala 401:37]
  wire [1:0] _GEN_125 = ocpSlaveReg_Resp == 2'h3 ? _T_10 : _GEN_112; // @[MCache.scala 451:43 MCache.scala 454:17]
  wire [2:0] _GEN_126 = ocpSlaveReg_Resp == 2'h3 ? 3'h3 : _GEN_119; // @[MCache.scala 451:43 MCache.scala 455:14]
  wire [2:0] _GEN_129 = _T_16 ? 3'h4 : _GEN_126; // @[MCache.scala 462:51 MCache.scala 465:16]
  wire  _GEN_131 = stateReg == 3'h3 & _T_16; // @[MCache.scala 458:34 MCache.scala 449:13]
  wire [2:0] _GEN_132 = stateReg == 3'h3 ? _GEN_129 : _GEN_126; // @[MCache.scala 458:34]
  wire  _GEN_133 = stateReg == 3'h4 | _GEN_131; // @[MCache.scala 469:37 MCache.scala 470:19]
  wire  _GEN_135 = stateReg == 3'h5 | _GEN_133; // @[MCache.scala 473:37 MCache.scala 474:19]
  wire [31:0] callRetBaseNext = io_exmcache_doCallRet ? io_exmcache_callRetBase : callRetBaseReg; // @[MCache.scala 341:32 MCache.scala 342:21 MCache.scala 326:19]
  assign io_fetchEna = stateReg == 3'h2 ? _GEN_103 : _GEN_49; // @[MCache.scala 401:37]
  assign io_ctrlrepl_wEna = stateReg == 3'h2 & _GEN_108; // @[MCache.scala 401:37 MCache.scala 322:8]
  assign io_ctrlrepl_wData = stateReg == 3'h2 ? _GEN_107 : {{20'd0}, _GEN_58}; // @[MCache.scala 401:37]
  assign io_ctrlrepl_wAddr = stateReg == 3'h2 ? _GEN_109 : _GEN_59; // @[MCache.scala 401:37]
  assign io_ctrlrepl_wTag = stateReg == 3'h1 & _GEN_45; // @[MCache.scala 371:33 MCache.scala 321:8]
  assign io_ctrlrepl_addrEven = addrEven[10:0]; // @[MCache.scala 483:24]
  assign io_ctrlrepl_addrOdd = addrOdd[10:0]; // @[MCache.scala 484:23]
  assign io_ctrlrepl_instrStall = stateReg != 3'h0; // @[MCache.scala 489:38]
  assign io_ocp_port_M_Cmd = ocpSlaveReg_Resp == 2'h3 ? 3'h0 : _GEN_113; // @[MCache.scala 451:43 MCache.scala 452:23]
  assign io_ocp_port_M_Addr = _GEN_115[31:0];
  assign io_illMem = stateReg == 3'h3 & _T_16; // @[MCache.scala 458:34 MCache.scala 449:13]
  assign io_forceHit = stateReg == 3'h6 | _GEN_135; // @[MCache.scala 477:37 MCache.scala 478:19]
  always @(posedge clock) begin
    if (reset) begin // @[MCache.scala 293:21]
      stateReg <= 3'h0; // @[MCache.scala 293:21]
    end else if (stateReg == 3'h6) begin // @[MCache.scala 477:37]
      stateReg <= 3'h0; // @[MCache.scala 479:16]
    end else if (stateReg == 3'h5) begin // @[MCache.scala 473:37]
      stateReg <= 3'h6; // @[MCache.scala 475:16]
    end else if (stateReg == 3'h4) begin // @[MCache.scala 469:37]
      stateReg <= 3'h5; // @[MCache.scala 471:16]
    end else begin
      stateReg <= _GEN_132;
    end
    if (reset) begin // @[MCache.scala 302:22]
      ocpCmdReg <= 3'h0; // @[MCache.scala 302:22]
    end else if (ocpSlaveReg_Resp == 2'h3) begin // @[MCache.scala 451:43]
      ocpCmdReg <= 3'h0; // @[MCache.scala 453:15]
    end else if (stateReg == 3'h2) begin // @[MCache.scala 401:37]
      if (fetchCntReg <= transferSizeReg) begin // @[MCache.scala 403:43]
        ocpCmdReg <= _GEN_83;
      end else begin
        ocpCmdReg <= _GEN_54;
      end
    end else begin
      ocpCmdReg <= _GEN_54;
    end
    if (stateReg == 3'h2) begin // @[MCache.scala 401:37]
      if (fetchCntReg <= transferSizeReg) begin // @[MCache.scala 403:43]
        if (_T_8) begin // @[MCache.scala 404:47]
          if (fetchCntReg < transferSizeReg) begin // @[MCache.scala 407:45]
            ocpAddrReg <= _GEN_65;
          end else begin
            ocpAddrReg <= _GEN_56;
          end
        end else begin
          ocpAddrReg <= _GEN_56;
        end
      end else begin
        ocpAddrReg <= _GEN_56;
      end
    end else begin
      ocpAddrReg <= _GEN_56;
    end
    transferSizeReg <= _GEN_51[10:0];
    if (stateReg == 3'h2) begin // @[MCache.scala 401:37]
      if (fetchCntReg <= transferSizeReg) begin // @[MCache.scala 403:43]
        if (_T_8) begin // @[MCache.scala 404:47]
          fetchCntReg <= _T_26; // @[MCache.scala 405:21]
        end else begin
          fetchCntReg <= _GEN_52;
        end
      end else begin
        fetchCntReg <= _GEN_52;
      end
    end else begin
      fetchCntReg <= _GEN_52;
    end
    if (stateReg == 3'h3) begin // @[MCache.scala 458:34]
      if (ocpSlaveReg_Resp != 2'h0) begin // @[MCache.scala 459:46]
        burstCntReg <= _T_10; // @[MCache.scala 460:19]
      end else begin
        burstCntReg <= _GEN_125;
      end
    end else begin
      burstCntReg <= _GEN_125;
    end
    callRetBaseReg <= callRetBaseNext; // @[MCache.scala 327:18]
    if (io_exmcache_doCallRet) begin // @[MCache.scala 341:32]
      addrEvenReg <= io_femcache_addrEven; // @[MCache.scala 343:17]
    end
    if (io_exmcache_doCallRet) begin // @[MCache.scala 341:32]
      addrOddReg <= io_femcache_addrOdd; // @[MCache.scala 344:16]
    end
    ocpSlaveReg_Resp <= io_ocp_port_S_Resp; // @[MCache.scala 315:24]
    ocpSlaveReg_Data <= io_ocp_port_S_Data; // @[MCache.scala 315:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  ocpCmdReg = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  ocpAddrReg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  transferSizeReg = _RAND_3[10:0];
  _RAND_4 = {1{`RANDOM}};
  fetchCntReg = _RAND_4[10:0];
  _RAND_5 = {1{`RANDOM}};
  burstCntReg = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  callRetBaseReg = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  addrEvenReg = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  addrOddReg = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  ocpSlaveReg_Resp = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  ocpSlaveReg_Data = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MCacheReplFifo(
  input         clock,
  input         reset,
  input         io_ena_in,
  input         io_invalidate,
  output        io_hitEna,
  input         io_exmcache_doCallRet,
  input  [31:0] io_exmcache_callRetBase,
  input  [31:0] io_exmcache_callRetAddr,
  output [31:0] io_mcachefe_instrEven,
  output [31:0] io_mcachefe_instrOdd,
  output [31:0] io_mcachefe_base,
  output [10:0] io_mcachefe_relBase,
  output [11:0] io_mcachefe_relPc,
  output [31:0] io_mcachefe_reloc,
  output [1:0]  io_mcachefe_memSel,
  input         io_ctrlrepl_wEna,
  input  [31:0] io_ctrlrepl_wData,
  input  [31:0] io_ctrlrepl_wAddr,
  input         io_ctrlrepl_wTag,
  input  [10:0] io_ctrlrepl_addrEven,
  input  [10:0] io_ctrlrepl_addrOdd,
  input         io_ctrlrepl_instrStall,
  output        io_replctrl_hit,
  output        io_memIn_wEven,
  output        io_memIn_wOdd,
  output [31:0] io_memIn_wData,
  output [9:0]  io_memIn_wAddr,
  output [9:0]  io_memIn_addrEven,
  output [9:0]  io_memIn_addrOdd,
  input  [31:0] io_memOut_instrEven,
  input  [31:0] io_memOut_instrOdd
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] nextIndexReg; // @[MCache.scala 146:25]
  reg [3:0] nextTagReg; // @[MCache.scala 147:23]
  reg [10:0] nextPosReg; // @[MCache.scala 148:23]
  reg [12:0] freeSpaceReg; // @[MCache.scala 149:25]
  reg [10:0] posReg; // @[MCache.scala 151:19]
  reg  hitReg; // @[MCache.scala 152:19]
  reg [10:0] wrPosReg; // @[MCache.scala 154:21]
  reg [31:0] callRetBaseReg; // @[MCache.scala 155:27]
  reg [31:0] callAddrReg; // @[MCache.scala 157:24]
  reg  selSpmReg; // @[MCache.scala 158:22]
  reg  selCacheReg; // @[MCache.scala 160:24]
  wire [31:0] _GEN_94 = 4'h0 == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_0 = io_ctrlrepl_wTag ? _GEN_94 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_110 = 4'h0 == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_178 = io_ctrlrepl_wTag & _GEN_110; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_229 = 4'h0 == nextTagReg ? 1'h0 : _GEN_178; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_262 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_229 : _GEN_178; // @[MCache.scala 238:33]
  wire  validVec_0 = io_invalidate ? 1'h0 : _GEN_262; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_0 = io_exmcache_callRetBase == addrVec_0 & validVec_0; // @[MCache.scala 179:50]
  wire [10:0] _GEN_62 = 4'h0 == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_0 = io_ctrlrepl_wTag ? _GEN_62 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_0 = hitVec_0 ? posVec_0 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_95 = 4'h1 == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_1 = io_ctrlrepl_wTag ? _GEN_95 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_111 = 4'h1 == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_179 = io_ctrlrepl_wTag & _GEN_111; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_230 = 4'h1 == nextTagReg ? 1'h0 : _GEN_179; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_263 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_230 : _GEN_179; // @[MCache.scala 238:33]
  wire  validVec_1 = io_invalidate ? 1'h0 : _GEN_263; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_1 = io_exmcache_callRetBase == addrVec_1 & validVec_1; // @[MCache.scala 179:50]
  wire [10:0] _GEN_63 = 4'h1 == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_1 = io_ctrlrepl_wTag ? _GEN_63 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_1 = hitVec_1 ? posVec_1 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_96 = 4'h2 == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_2 = io_ctrlrepl_wTag ? _GEN_96 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_112 = 4'h2 == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_180 = io_ctrlrepl_wTag & _GEN_112; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_231 = 4'h2 == nextTagReg ? 1'h0 : _GEN_180; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_264 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_231 : _GEN_180; // @[MCache.scala 238:33]
  wire  validVec_2 = io_invalidate ? 1'h0 : _GEN_264; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_2 = io_exmcache_callRetBase == addrVec_2 & validVec_2; // @[MCache.scala 179:50]
  wire [10:0] _GEN_64 = 4'h2 == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_2 = io_ctrlrepl_wTag ? _GEN_64 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_2 = hitVec_2 ? posVec_2 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_97 = 4'h3 == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_3 = io_ctrlrepl_wTag ? _GEN_97 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_113 = 4'h3 == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_181 = io_ctrlrepl_wTag & _GEN_113; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_232 = 4'h3 == nextTagReg ? 1'h0 : _GEN_181; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_265 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_232 : _GEN_181; // @[MCache.scala 238:33]
  wire  validVec_3 = io_invalidate ? 1'h0 : _GEN_265; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_3 = io_exmcache_callRetBase == addrVec_3 & validVec_3; // @[MCache.scala 179:50]
  wire [10:0] _GEN_65 = 4'h3 == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_3 = io_ctrlrepl_wTag ? _GEN_65 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_3 = hitVec_3 ? posVec_3 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_98 = 4'h4 == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_4 = io_ctrlrepl_wTag ? _GEN_98 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_114 = 4'h4 == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_182 = io_ctrlrepl_wTag & _GEN_114; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_233 = 4'h4 == nextTagReg ? 1'h0 : _GEN_182; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_266 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_233 : _GEN_182; // @[MCache.scala 238:33]
  wire  validVec_4 = io_invalidate ? 1'h0 : _GEN_266; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_4 = io_exmcache_callRetBase == addrVec_4 & validVec_4; // @[MCache.scala 179:50]
  wire [10:0] _GEN_66 = 4'h4 == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_4 = io_ctrlrepl_wTag ? _GEN_66 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_4 = hitVec_4 ? posVec_4 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_99 = 4'h5 == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_5 = io_ctrlrepl_wTag ? _GEN_99 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_115 = 4'h5 == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_183 = io_ctrlrepl_wTag & _GEN_115; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_234 = 4'h5 == nextTagReg ? 1'h0 : _GEN_183; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_267 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_234 : _GEN_183; // @[MCache.scala 238:33]
  wire  validVec_5 = io_invalidate ? 1'h0 : _GEN_267; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_5 = io_exmcache_callRetBase == addrVec_5 & validVec_5; // @[MCache.scala 179:50]
  wire [10:0] _GEN_67 = 4'h5 == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_5 = io_ctrlrepl_wTag ? _GEN_67 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_5 = hitVec_5 ? posVec_5 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_100 = 4'h6 == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_6 = io_ctrlrepl_wTag ? _GEN_100 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_116 = 4'h6 == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_184 = io_ctrlrepl_wTag & _GEN_116; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_235 = 4'h6 == nextTagReg ? 1'h0 : _GEN_184; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_268 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_235 : _GEN_184; // @[MCache.scala 238:33]
  wire  validVec_6 = io_invalidate ? 1'h0 : _GEN_268; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_6 = io_exmcache_callRetBase == addrVec_6 & validVec_6; // @[MCache.scala 179:50]
  wire [10:0] _GEN_68 = 4'h6 == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_6 = io_ctrlrepl_wTag ? _GEN_68 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_6 = hitVec_6 ? posVec_6 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_101 = 4'h7 == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_7 = io_ctrlrepl_wTag ? _GEN_101 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_117 = 4'h7 == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_185 = io_ctrlrepl_wTag & _GEN_117; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_236 = 4'h7 == nextTagReg ? 1'h0 : _GEN_185; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_269 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_236 : _GEN_185; // @[MCache.scala 238:33]
  wire  validVec_7 = io_invalidate ? 1'h0 : _GEN_269; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_7 = io_exmcache_callRetBase == addrVec_7 & validVec_7; // @[MCache.scala 179:50]
  wire [10:0] _GEN_69 = 4'h7 == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_7 = io_ctrlrepl_wTag ? _GEN_69 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_7 = hitVec_7 ? posVec_7 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_102 = 4'h8 == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_8 = io_ctrlrepl_wTag ? _GEN_102 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_118 = 4'h8 == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_186 = io_ctrlrepl_wTag & _GEN_118; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_237 = 4'h8 == nextTagReg ? 1'h0 : _GEN_186; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_270 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_237 : _GEN_186; // @[MCache.scala 238:33]
  wire  validVec_8 = io_invalidate ? 1'h0 : _GEN_270; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_8 = io_exmcache_callRetBase == addrVec_8 & validVec_8; // @[MCache.scala 179:50]
  wire [10:0] _GEN_70 = 4'h8 == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_8 = io_ctrlrepl_wTag ? _GEN_70 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_8 = hitVec_8 ? posVec_8 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_103 = 4'h9 == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_9 = io_ctrlrepl_wTag ? _GEN_103 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_119 = 4'h9 == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_187 = io_ctrlrepl_wTag & _GEN_119; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_238 = 4'h9 == nextTagReg ? 1'h0 : _GEN_187; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_271 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_238 : _GEN_187; // @[MCache.scala 238:33]
  wire  validVec_9 = io_invalidate ? 1'h0 : _GEN_271; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_9 = io_exmcache_callRetBase == addrVec_9 & validVec_9; // @[MCache.scala 179:50]
  wire [10:0] _GEN_71 = 4'h9 == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_9 = io_ctrlrepl_wTag ? _GEN_71 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_9 = hitVec_9 ? posVec_9 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_104 = 4'ha == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_10 = io_ctrlrepl_wTag ? _GEN_104 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_120 = 4'ha == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_188 = io_ctrlrepl_wTag & _GEN_120; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_239 = 4'ha == nextTagReg ? 1'h0 : _GEN_188; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_272 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_239 : _GEN_188; // @[MCache.scala 238:33]
  wire  validVec_10 = io_invalidate ? 1'h0 : _GEN_272; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_10 = io_exmcache_callRetBase == addrVec_10 & validVec_10; // @[MCache.scala 179:50]
  wire [10:0] _GEN_72 = 4'ha == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_10 = io_ctrlrepl_wTag ? _GEN_72 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_10 = hitVec_10 ? posVec_10 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_105 = 4'hb == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_11 = io_ctrlrepl_wTag ? _GEN_105 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_121 = 4'hb == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_189 = io_ctrlrepl_wTag & _GEN_121; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_240 = 4'hb == nextTagReg ? 1'h0 : _GEN_189; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_273 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_240 : _GEN_189; // @[MCache.scala 238:33]
  wire  validVec_11 = io_invalidate ? 1'h0 : _GEN_273; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_11 = io_exmcache_callRetBase == addrVec_11 & validVec_11; // @[MCache.scala 179:50]
  wire [10:0] _GEN_73 = 4'hb == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_11 = io_ctrlrepl_wTag ? _GEN_73 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_11 = hitVec_11 ? posVec_11 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_106 = 4'hc == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_12 = io_ctrlrepl_wTag ? _GEN_106 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_122 = 4'hc == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_190 = io_ctrlrepl_wTag & _GEN_122; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_241 = 4'hc == nextTagReg ? 1'h0 : _GEN_190; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_274 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_241 : _GEN_190; // @[MCache.scala 238:33]
  wire  validVec_12 = io_invalidate ? 1'h0 : _GEN_274; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_12 = io_exmcache_callRetBase == addrVec_12 & validVec_12; // @[MCache.scala 179:50]
  wire [10:0] _GEN_74 = 4'hc == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_12 = io_ctrlrepl_wTag ? _GEN_74 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_12 = hitVec_12 ? posVec_12 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_107 = 4'hd == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_13 = io_ctrlrepl_wTag ? _GEN_107 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_123 = 4'hd == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_191 = io_ctrlrepl_wTag & _GEN_123; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_242 = 4'hd == nextTagReg ? 1'h0 : _GEN_191; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_275 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_242 : _GEN_191; // @[MCache.scala 238:33]
  wire  validVec_13 = io_invalidate ? 1'h0 : _GEN_275; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_13 = io_exmcache_callRetBase == addrVec_13 & validVec_13; // @[MCache.scala 179:50]
  wire [10:0] _GEN_75 = 4'hd == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_13 = io_ctrlrepl_wTag ? _GEN_75 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_13 = hitVec_13 ? posVec_13 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_108 = 4'he == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_14 = io_ctrlrepl_wTag ? _GEN_108 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_124 = 4'he == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_192 = io_ctrlrepl_wTag & _GEN_124; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_243 = 4'he == nextTagReg ? 1'h0 : _GEN_192; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_276 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_243 : _GEN_192; // @[MCache.scala 238:33]
  wire  validVec_14 = io_invalidate ? 1'h0 : _GEN_276; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_14 = io_exmcache_callRetBase == addrVec_14 & validVec_14; // @[MCache.scala 179:50]
  wire [10:0] _GEN_76 = 4'he == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_14 = io_ctrlrepl_wTag ? _GEN_76 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_14 = hitVec_14 ? posVec_14 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire [31:0] _GEN_109 = 4'hf == nextIndexReg ? io_ctrlrepl_wAddr : 32'h0; // @[MCache.scala 227:27 MCache.scala 227:27 compatibility.scala 127:12]
  wire [31:0] addrVec_15 = io_ctrlrepl_wTag ? _GEN_109 : 32'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_125 = 4'hf == nextIndexReg; // @[MCache.scala 228:28 MCache.scala 228:28 compatibility.scala 127:12]
  wire  _GEN_193 = io_ctrlrepl_wTag & _GEN_125; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire  _GEN_244 = 4'hf == nextTagReg ? 1'h0 : _GEN_193; // @[MCache.scala 241:26 MCache.scala 241:26]
  wire  _GEN_277 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_244 : _GEN_193; // @[MCache.scala 238:33]
  wire  validVec_15 = io_invalidate ? 1'h0 : _GEN_277; // @[MCache.scala 279:24 MCache.scala 280:20]
  wire  hitVec_15 = io_exmcache_callRetBase == addrVec_15 & validVec_15; // @[MCache.scala 179:50]
  wire [10:0] _GEN_77 = 4'hf == nextIndexReg ? nextPosReg : 11'h0; // @[MCache.scala 225:26 MCache.scala 225:26 compatibility.scala 127:12]
  wire [10:0] posVec_15 = io_ctrlrepl_wTag ? _GEN_77 : 11'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [10:0] mergePosVec_15 = hitVec_15 ? posVec_15 : 11'h0; // @[MCache.scala 179:66 MCache.scala 181:22 MCache.scala 178:20]
  wire  hit = hitVec_0 | hitVec_1 | hitVec_2 | hitVec_3 | hitVec_4 | hitVec_5 | hitVec_6 | hitVec_7 | hitVec_8 |
    hitVec_9 | hitVec_10 | hitVec_11 | hitVec_12 | hitVec_13 | hitVec_14 | hitVec_15; // @[MCache.scala 184:39]
  wire [10:0] _T_48 = mergePosVec_0 | mergePosVec_1; // @[MCache.scala 185:49]
  wire [10:0] _T_49 = _T_48 | mergePosVec_2; // @[MCache.scala 185:49]
  wire [10:0] _T_50 = _T_49 | mergePosVec_3; // @[MCache.scala 185:49]
  wire [10:0] _T_51 = _T_50 | mergePosVec_4; // @[MCache.scala 185:49]
  wire [10:0] _T_52 = _T_51 | mergePosVec_5; // @[MCache.scala 185:49]
  wire [10:0] _T_53 = _T_52 | mergePosVec_6; // @[MCache.scala 185:49]
  wire [10:0] _T_54 = _T_53 | mergePosVec_7; // @[MCache.scala 185:49]
  wire [10:0] _T_55 = _T_54 | mergePosVec_8; // @[MCache.scala 185:49]
  wire [10:0] _T_56 = _T_55 | mergePosVec_9; // @[MCache.scala 185:49]
  wire [10:0] _T_57 = _T_56 | mergePosVec_10; // @[MCache.scala 185:49]
  wire [10:0] _T_58 = _T_57 | mergePosVec_11; // @[MCache.scala 185:49]
  wire [10:0] _T_59 = _T_58 | mergePosVec_12; // @[MCache.scala 185:49]
  wire [10:0] _T_60 = _T_59 | mergePosVec_13; // @[MCache.scala 185:49]
  wire [10:0] _T_61 = _T_60 | mergePosVec_14; // @[MCache.scala 185:49]
  wire [10:0] _T_62 = _T_61 | mergePosVec_15; // @[MCache.scala 185:49]
  wire  _T_67 = io_exmcache_callRetBase[31:15] >= 17'h1; // @[MCache.scala 193:74]
  wire  _GEN_34 = _T_67 ? hit : hitReg; // @[MCache.scala 195:21 MCache.scala 196:15 MCache.scala 165:11]
  wire  _GEN_42 = io_exmcache_doCallRet & io_ena_in ? _GEN_34 : hitReg; // @[MCache.scala 188:45 MCache.scala 165:11]
  wire [13:0] relBase = selCacheReg ? {{3'd0}, posReg} : callRetBaseReg[13:0]; // @[MCache.scala 207:20]
  wire [31:0] _GEN_297 = {{18'd0}, relBase}; // @[MCache.scala 210:27]
  wire [31:0] relPc = callAddrReg + _GEN_297; // @[MCache.scala 210:27]
  wire [31:0] _GEN_298 = {{21'd0}, posReg}; // @[MCache.scala 213:34]
  wire [31:0] _T_71 = callRetBaseReg - _GEN_298; // @[MCache.scala 213:34]
  wire [14:0] _T_72 = selSpmReg ? 15'h4000 : 15'h0; // @[MCache.scala 214:22]
  wire [11:0] _T_74 = io_ctrlrepl_wData[11:0]; // @[MCache.scala 223:75]
  wire [12:0] _GEN_299 = {{1{_T_74[11]}},_T_74}; // @[MCache.scala 223:34]
  wire [12:0] _T_77 = $signed(freeSpaceReg) - $signed(_GEN_299); // @[MCache.scala 223:34]
  wire [11:0] _GEN_78 = 4'h0 == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_146 = io_ctrlrepl_wTag ? _GEN_78 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_213 = 4'h0 == nextTagReg ? 12'h0 : _GEN_146; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_0 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_213 : _GEN_146; // @[MCache.scala 238:33]
  wire [11:0] _GEN_79 = 4'h1 == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_147 = io_ctrlrepl_wTag ? _GEN_79 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_214 = 4'h1 == nextTagReg ? 12'h0 : _GEN_147; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_1 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_214 : _GEN_147; // @[MCache.scala 238:33]
  wire [11:0] _GEN_47 = 4'h1 == nextIndexReg ? sizeVec_1 : sizeVec_0; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_80 = 4'h2 == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_148 = io_ctrlrepl_wTag ? _GEN_80 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_215 = 4'h2 == nextTagReg ? 12'h0 : _GEN_148; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_2 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_215 : _GEN_148; // @[MCache.scala 238:33]
  wire [11:0] _GEN_48 = 4'h2 == nextIndexReg ? sizeVec_2 : _GEN_47; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_81 = 4'h3 == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_149 = io_ctrlrepl_wTag ? _GEN_81 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_216 = 4'h3 == nextTagReg ? 12'h0 : _GEN_149; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_3 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_216 : _GEN_149; // @[MCache.scala 238:33]
  wire [11:0] _GEN_49 = 4'h3 == nextIndexReg ? sizeVec_3 : _GEN_48; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_82 = 4'h4 == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_150 = io_ctrlrepl_wTag ? _GEN_82 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_217 = 4'h4 == nextTagReg ? 12'h0 : _GEN_150; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_4 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_217 : _GEN_150; // @[MCache.scala 238:33]
  wire [11:0] _GEN_50 = 4'h4 == nextIndexReg ? sizeVec_4 : _GEN_49; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_83 = 4'h5 == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_151 = io_ctrlrepl_wTag ? _GEN_83 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_218 = 4'h5 == nextTagReg ? 12'h0 : _GEN_151; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_5 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_218 : _GEN_151; // @[MCache.scala 238:33]
  wire [11:0] _GEN_51 = 4'h5 == nextIndexReg ? sizeVec_5 : _GEN_50; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_84 = 4'h6 == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_152 = io_ctrlrepl_wTag ? _GEN_84 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_219 = 4'h6 == nextTagReg ? 12'h0 : _GEN_152; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_6 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_219 : _GEN_152; // @[MCache.scala 238:33]
  wire [11:0] _GEN_52 = 4'h6 == nextIndexReg ? sizeVec_6 : _GEN_51; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_85 = 4'h7 == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_153 = io_ctrlrepl_wTag ? _GEN_85 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_220 = 4'h7 == nextTagReg ? 12'h0 : _GEN_153; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_7 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_220 : _GEN_153; // @[MCache.scala 238:33]
  wire [11:0] _GEN_53 = 4'h7 == nextIndexReg ? sizeVec_7 : _GEN_52; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_86 = 4'h8 == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_154 = io_ctrlrepl_wTag ? _GEN_86 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_221 = 4'h8 == nextTagReg ? 12'h0 : _GEN_154; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_8 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_221 : _GEN_154; // @[MCache.scala 238:33]
  wire [11:0] _GEN_54 = 4'h8 == nextIndexReg ? sizeVec_8 : _GEN_53; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_87 = 4'h9 == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_155 = io_ctrlrepl_wTag ? _GEN_87 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_222 = 4'h9 == nextTagReg ? 12'h0 : _GEN_155; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_9 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_222 : _GEN_155; // @[MCache.scala 238:33]
  wire [11:0] _GEN_55 = 4'h9 == nextIndexReg ? sizeVec_9 : _GEN_54; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_88 = 4'ha == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_156 = io_ctrlrepl_wTag ? _GEN_88 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_223 = 4'ha == nextTagReg ? 12'h0 : _GEN_156; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_10 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_223 : _GEN_156; // @[MCache.scala 238:33]
  wire [11:0] _GEN_56 = 4'ha == nextIndexReg ? sizeVec_10 : _GEN_55; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_89 = 4'hb == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_157 = io_ctrlrepl_wTag ? _GEN_89 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_224 = 4'hb == nextTagReg ? 12'h0 : _GEN_157; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_11 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_224 : _GEN_157; // @[MCache.scala 238:33]
  wire [11:0] _GEN_57 = 4'hb == nextIndexReg ? sizeVec_11 : _GEN_56; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_90 = 4'hc == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_158 = io_ctrlrepl_wTag ? _GEN_90 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_225 = 4'hc == nextTagReg ? 12'h0 : _GEN_158; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_12 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_225 : _GEN_158; // @[MCache.scala 238:33]
  wire [11:0] _GEN_58 = 4'hc == nextIndexReg ? sizeVec_12 : _GEN_57; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_91 = 4'hd == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_159 = io_ctrlrepl_wTag ? _GEN_91 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_226 = 4'hd == nextTagReg ? 12'h0 : _GEN_159; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_13 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_226 : _GEN_159; // @[MCache.scala 238:33]
  wire [11:0] _GEN_59 = 4'hd == nextIndexReg ? sizeVec_13 : _GEN_58; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_92 = 4'he == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_160 = io_ctrlrepl_wTag ? _GEN_92 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_227 = 4'he == nextTagReg ? 12'h0 : _GEN_160; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_14 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_227 : _GEN_160; // @[MCache.scala 238:33]
  wire [11:0] _GEN_60 = 4'he == nextIndexReg ? sizeVec_14 : _GEN_59; // @[MCache.scala 223:106 MCache.scala 223:106]
  wire [11:0] _GEN_93 = 4'hf == nextIndexReg ? io_ctrlrepl_wData[11:0] : 12'h0; // @[MCache.scala 226:27 MCache.scala 226:27 compatibility.scala 127:12]
  wire [11:0] _GEN_161 = io_ctrlrepl_wTag ? _GEN_93 : 12'h0; // @[MCache.scala 219:27 compatibility.scala 127:12]
  wire [11:0] _GEN_228 = 4'hf == nextTagReg ? 12'h0 : _GEN_161; // @[MCache.scala 240:25 MCache.scala 240:25]
  wire [11:0] sizeVec_15 = $signed(freeSpaceReg) < 13'sh0 ? _GEN_228 : _GEN_161; // @[MCache.scala 238:33]
  wire [11:0] _T_78 = 4'hf == nextIndexReg ? sizeVec_15 : _GEN_60; // @[MCache.scala 223:106]
  wire [12:0] _GEN_300 = {{1{_T_78[11]}},_T_78}; // @[MCache.scala 223:82]
  wire [12:0] _T_81 = $signed(_T_77) + $signed(_GEN_300); // @[MCache.scala 223:82]
  wire [10:0] _T_85 = nextPosReg + io_ctrlrepl_wData[10:0]; // @[MCache.scala 230:30]
  wire [3:0] _T_88 = nextIndexReg + 4'h1; // @[MCache.scala 231:86]
  wire [3:0] _T_89 = nextIndexReg == 4'hf ? 4'h0 : _T_88; // @[MCache.scala 231:22]
  wire [11:0] _GEN_198 = 4'h1 == nextTagReg ? sizeVec_1 : sizeVec_0; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_199 = 4'h2 == nextTagReg ? sizeVec_2 : _GEN_198; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_200 = 4'h3 == nextTagReg ? sizeVec_3 : _GEN_199; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_201 = 4'h4 == nextTagReg ? sizeVec_4 : _GEN_200; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_202 = 4'h5 == nextTagReg ? sizeVec_5 : _GEN_201; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_203 = 4'h6 == nextTagReg ? sizeVec_6 : _GEN_202; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_204 = 4'h7 == nextTagReg ? sizeVec_7 : _GEN_203; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_205 = 4'h8 == nextTagReg ? sizeVec_8 : _GEN_204; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_206 = 4'h9 == nextTagReg ? sizeVec_9 : _GEN_205; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_207 = 4'ha == nextTagReg ? sizeVec_10 : _GEN_206; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_208 = 4'hb == nextTagReg ? sizeVec_11 : _GEN_207; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_209 = 4'hc == nextTagReg ? sizeVec_12 : _GEN_208; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_210 = 4'hd == nextTagReg ? sizeVec_13 : _GEN_209; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _GEN_211 = 4'he == nextTagReg ? sizeVec_14 : _GEN_210; // @[MCache.scala 239:56 MCache.scala 239:56]
  wire [11:0] _T_92 = 4'hf == nextTagReg ? sizeVec_15 : _GEN_211; // @[MCache.scala 239:56]
  wire [12:0] _GEN_301 = {{1{_T_92[11]}},_T_92}; // @[MCache.scala 239:34]
  wire [12:0] _T_95 = $signed(freeSpaceReg) + $signed(_GEN_301); // @[MCache.scala 239:34]
  wire [3:0] _T_98 = nextTagReg + 4'h1; // @[MCache.scala 242:82]
  wire  wParity = io_ctrlrepl_wAddr[0]; // @[MCache.scala 245:34]
  wire [31:0] _GEN_302 = {{21'd0}, wrPosReg}; // @[MCache.scala 247:25]
  wire [31:0] _T_101 = _GEN_302 + io_ctrlrepl_wAddr; // @[MCache.scala 247:25]
  reg [31:0] instrEvenReg; // @[MCache.scala 258:25]
  reg [31:0] instrOddReg; // @[MCache.scala 259:24]
  wire  hitNext = io_ctrlrepl_wTag | _GEN_42; // @[MCache.scala 219:27 MCache.scala 220:13]
  wire [31:0] callRetBaseNext = io_exmcache_doCallRet & io_ena_in ? io_exmcache_callRetBase : callRetBaseReg; // @[MCache.scala 188:45 MCache.scala 190:21 MCache.scala 167:19]
  wire  selSpmNext = io_exmcache_doCallRet & io_ena_in ? io_exmcache_callRetBase[31:14] == 18'h1 : selSpmReg; // @[MCache.scala 188:45 MCache.scala 192:16 MCache.scala 169:14]
  wire  selCacheNext = io_exmcache_doCallRet & io_ena_in ? _T_67 : selCacheReg; // @[MCache.scala 188:45 MCache.scala 194:18 MCache.scala 171:16]
  assign io_hitEna = hitReg; // @[MCache.scala 276:13]
  assign io_mcachefe_instrEven = io_ctrlrepl_instrStall ? instrEvenReg : io_memOut_instrEven; // @[MCache.scala 266:31]
  assign io_mcachefe_instrOdd = io_ctrlrepl_instrStall ? instrOddReg : io_memOut_instrOdd; // @[MCache.scala 267:30]
  assign io_mcachefe_base = callRetBaseReg; // @[MCache.scala 268:20]
  assign io_mcachefe_relBase = relBase[10:0]; // @[MCache.scala 269:23]
  assign io_mcachefe_relPc = relPc[11:0]; // @[MCache.scala 270:21]
  assign io_mcachefe_reloc = selCacheReg ? _T_71 : {{17'd0}, _T_72}; // @[MCache.scala 212:18]
  assign io_mcachefe_memSel = {selSpmReg,selCacheReg}; // @[Cat.scala 30:58]
  assign io_replctrl_hit = hitReg; // @[MCache.scala 274:19]
  assign io_memIn_wEven = wParity ? 1'h0 : io_ctrlrepl_wEna; // @[MCache.scala 251:24]
  assign io_memIn_wOdd = wParity & io_ctrlrepl_wEna; // @[MCache.scala 252:23]
  assign io_memIn_wData = io_ctrlrepl_wData; // @[MCache.scala 253:18]
  assign io_memIn_wAddr = _T_101[10:1]; // @[MCache.scala 247:45]
  assign io_memIn_addrEven = io_ctrlrepl_addrEven[10:1]; // @[MCache.scala 248:40]
  assign io_memIn_addrOdd = io_ctrlrepl_addrOdd[10:1]; // @[MCache.scala 249:38]
  always @(posedge clock) begin
    if (reset) begin // @[MCache.scala 146:25]
      nextIndexReg <= 4'h0; // @[MCache.scala 146:25]
    end else if (io_ctrlrepl_wTag) begin // @[MCache.scala 219:27]
      if (nextIndexReg == 4'hf) begin // @[MCache.scala 231:22]
        nextIndexReg <= 4'h0;
      end else begin
        nextIndexReg <= _T_88;
      end
    end
    if (reset) begin // @[MCache.scala 147:23]
      nextTagReg <= 4'h0; // @[MCache.scala 147:23]
    end else if ($signed(freeSpaceReg) < 13'sh0) begin // @[MCache.scala 238:33]
      if (nextTagReg == 4'hf) begin // @[MCache.scala 242:22]
        nextTagReg <= 4'h0;
      end else begin
        nextTagReg <= _T_98;
      end
    end else if (io_ctrlrepl_wTag) begin // @[MCache.scala 219:27]
      if (nextTagReg == nextIndexReg) begin // @[MCache.scala 233:40]
        nextTagReg <= _T_89; // @[MCache.scala 234:18]
      end
    end
    if (reset) begin // @[MCache.scala 148:23]
      nextPosReg <= 11'h0; // @[MCache.scala 148:23]
    end else if (io_ctrlrepl_wTag) begin // @[MCache.scala 219:27]
      nextPosReg <= _T_85; // @[MCache.scala 230:16]
    end
    if (reset) begin // @[MCache.scala 149:25]
      freeSpaceReg <= 13'sh800; // @[MCache.scala 149:25]
    end else if ($signed(freeSpaceReg) < 13'sh0) begin // @[MCache.scala 238:33]
      freeSpaceReg <= _T_95; // @[MCache.scala 239:18]
    end else if (io_ctrlrepl_wTag) begin // @[MCache.scala 219:27]
      freeSpaceReg <= _T_81; // @[MCache.scala 223:18]
    end
    if (reset) begin // @[MCache.scala 151:19]
      posReg <= 11'h0; // @[MCache.scala 151:19]
    end else if (io_exmcache_doCallRet & io_ena_in) begin // @[MCache.scala 188:45]
      if (_T_67) begin // @[MCache.scala 195:21]
        if (hit) begin // @[MCache.scala 185:16]
          posReg <= _T_62;
        end else begin
          posReg <= nextPosReg;
        end
      end
    end
    hitReg <= reset | hitNext; // @[MCache.scala 152:19 MCache.scala 152:19 MCache.scala 166:10]
    if (reset) begin // @[MCache.scala 154:21]
      wrPosReg <= 11'h0; // @[MCache.scala 154:21]
    end else if (io_ctrlrepl_wTag) begin // @[MCache.scala 219:27]
      wrPosReg <= posReg; // @[MCache.scala 221:14]
    end
    if (reset) begin // @[MCache.scala 155:27]
      callRetBaseReg <= 32'h1; // @[MCache.scala 155:27]
    end else if (io_exmcache_doCallRet & io_ena_in) begin // @[MCache.scala 188:45]
      callRetBaseReg <= io_exmcache_callRetBase; // @[MCache.scala 190:21]
    end
    if (reset) begin // @[MCache.scala 157:24]
      callAddrReg <= 32'h1; // @[MCache.scala 157:24]
    end else if (io_exmcache_doCallRet & io_ena_in) begin // @[MCache.scala 188:45]
      callAddrReg <= io_exmcache_callRetAddr; // @[MCache.scala 191:17]
    end
    if (reset) begin // @[MCache.scala 158:22]
      selSpmReg <= 1'h0; // @[MCache.scala 158:22]
    end else if (io_exmcache_doCallRet & io_ena_in) begin // @[MCache.scala 188:45]
      selSpmReg <= io_exmcache_callRetBase[31:14] == 18'h1; // @[MCache.scala 192:16]
    end
    if (reset) begin // @[MCache.scala 160:24]
      selCacheReg <= 1'h0; // @[MCache.scala 160:24]
    end else if (io_exmcache_doCallRet & io_ena_in) begin // @[MCache.scala 188:45]
      selCacheReg <= _T_67; // @[MCache.scala 194:18]
    end
    if (~io_ctrlrepl_instrStall) begin // @[MCache.scala 262:34]
      instrEvenReg <= io_mcachefe_instrEven; // @[MCache.scala 263:18]
    end
    if (~io_ctrlrepl_instrStall) begin // @[MCache.scala 262:34]
      instrOddReg <= io_mcachefe_instrOdd; // @[MCache.scala 264:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  nextIndexReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  nextTagReg = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  nextPosReg = _RAND_2[10:0];
  _RAND_3 = {1{`RANDOM}};
  freeSpaceReg = _RAND_3[12:0];
  _RAND_4 = {1{`RANDOM}};
  posReg = _RAND_4[10:0];
  _RAND_5 = {1{`RANDOM}};
  hitReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  wrPosReg = _RAND_6[10:0];
  _RAND_7 = {1{`RANDOM}};
  callRetBaseReg = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  callAddrReg = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  selSpmReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  selCacheReg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  instrEvenReg = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  instrOddReg = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemBlock(
  input         clock,
  input  [9:0]  io_rdAddr,
  output [31:0] io_rdData,
  input  [9:0]  io_wrAddr,
  input         io_wrEna,
  input  [31:0] io_wrData
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:1023];
  wire [31:0] mem_MPORT_1_data;
  wire [9:0] mem_MPORT_1_addr;
  wire [31:0] mem_MPORT_data;
  wire [9:0] mem_MPORT_addr;
  wire  mem_MPORT_mask;
  wire  mem_MPORT_en;
  reg [9:0] rdAddrReg; // @[MemBlock.scala 59:22]
  reg  REG; // @[MemBlock.scala 64:14]
  reg [9:0] REG_1; // @[MemBlock.scala 65:14]
  wire  _T_4 = REG_1 == rdAddrReg; // @[MemBlock.scala 65:33]
  wire  _T_5 = REG & _T_4; // @[MemBlock.scala 64:44]
  reg [31:0] REG_2; // @[MemBlock.scala 66:29]
  assign mem_MPORT_1_addr = rdAddrReg;
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr];
  assign mem_MPORT_data = io_wrData;
  assign mem_MPORT_addr = io_wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEna;
  assign io_rdData = _T_5 ? REG_2 : mem_MPORT_1_data; // @[MemBlock.scala 65:48 MemBlock.scala 66:23 MemBlock.scala 60:13]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data;
    end
    rdAddrReg <= io_rdAddr; // @[MemBlock.scala 59:22]
    REG <= io_wrEna; // @[MemBlock.scala 64:14]
    REG_1 <= io_wrAddr; // @[MemBlock.scala 65:14]
    REG_2 <= io_wrData; // @[MemBlock.scala 66:29]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rdAddrReg = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_1 = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MCacheMem(
  input         clock,
  input         io_memIn_wEven,
  input         io_memIn_wOdd,
  input  [31:0] io_memIn_wData,
  input  [9:0]  io_memIn_wAddr,
  input  [9:0]  io_memIn_addrEven,
  input  [9:0]  io_memIn_addrOdd,
  output [31:0] io_memOut_instrEven,
  output [31:0] io_memOut_instrOdd
);
  wire  mcacheEven_clock; // @[MemBlock.scala 15:11]
  wire [9:0] mcacheEven_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [31:0] mcacheEven_io_rdData; // @[MemBlock.scala 15:11]
  wire [9:0] mcacheEven_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  mcacheEven_io_wrEna; // @[MemBlock.scala 15:11]
  wire [31:0] mcacheEven_io_wrData; // @[MemBlock.scala 15:11]
  wire  mcacheOdd_clock; // @[MemBlock.scala 15:11]
  wire [9:0] mcacheOdd_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [31:0] mcacheOdd_io_rdData; // @[MemBlock.scala 15:11]
  wire [9:0] mcacheOdd_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  mcacheOdd_io_wrEna; // @[MemBlock.scala 15:11]
  wire [31:0] mcacheOdd_io_wrData; // @[MemBlock.scala 15:11]
  MemBlock mcacheEven ( // @[MemBlock.scala 15:11]
    .clock(mcacheEven_clock),
    .io_rdAddr(mcacheEven_io_rdAddr),
    .io_rdData(mcacheEven_io_rdData),
    .io_wrAddr(mcacheEven_io_wrAddr),
    .io_wrEna(mcacheEven_io_wrEna),
    .io_wrData(mcacheEven_io_wrData)
  );
  MemBlock mcacheOdd ( // @[MemBlock.scala 15:11]
    .clock(mcacheOdd_clock),
    .io_rdAddr(mcacheOdd_io_rdAddr),
    .io_rdData(mcacheOdd_io_rdData),
    .io_wrAddr(mcacheOdd_io_wrAddr),
    .io_wrEna(mcacheOdd_io_wrEna),
    .io_wrData(mcacheOdd_io_wrData)
  );
  assign io_memOut_instrEven = mcacheEven_io_rdData; // @[MCache.scala 127:23]
  assign io_memOut_instrOdd = mcacheOdd_io_rdData; // @[MCache.scala 128:22]
  assign mcacheEven_clock = clock;
  assign mcacheEven_io_rdAddr = io_memIn_addrEven; // @[MemBlock.scala 44:12]
  assign mcacheEven_io_wrAddr = io_memIn_wAddr; // @[MemBlock.scala 34:12]
  assign mcacheEven_io_wrEna = io_memIn_wEven; // @[MemBlock.scala 35:11]
  assign mcacheEven_io_wrData = io_memIn_wData; // @[MemBlock.scala 36:12]
  assign mcacheOdd_clock = clock;
  assign mcacheOdd_io_rdAddr = io_memIn_addrOdd; // @[MemBlock.scala 44:12]
  assign mcacheOdd_io_wrAddr = io_memIn_wAddr; // @[MemBlock.scala 34:12]
  assign mcacheOdd_io_wrEna = io_memIn_wOdd; // @[MemBlock.scala 35:11]
  assign mcacheOdd_io_wrData = io_memIn_wData; // @[MemBlock.scala 36:12]
endmodule
module MCache(
  input         clock,
  input         reset,
  output        io_ena_out,
  input         io_ena_in,
  input         io_invalidate,
  input  [31:0] io_feicache_addrEven,
  input  [31:0] io_feicache_addrOdd,
  input         io_exicache_doCallRet,
  input  [31:0] io_exicache_callRetBase,
  input  [31:0] io_exicache_callRetAddr,
  output [31:0] io_icachefe_instrEven,
  output [31:0] io_icachefe_instrOdd,
  output [31:0] io_icachefe_base,
  output [10:0] io_icachefe_relBase,
  output [11:0] io_icachefe_relPc,
  output [31:0] io_icachefe_reloc,
  output [1:0]  io_icachefe_memSel,
  output [2:0]  io_ocp_port_M_Cmd,
  output [31:0] io_ocp_port_M_Addr,
  input  [1:0]  io_ocp_port_S_Resp,
  input  [31:0] io_ocp_port_S_Data,
  input         io_ocp_port_S_CmdAccept,
  output        io_illMem
);
  wire  ctrl_clock; // @[MCache.scala 86:20]
  wire  ctrl_reset; // @[MCache.scala 86:20]
  wire  ctrl_io_fetchEna; // @[MCache.scala 86:20]
  wire  ctrl_io_ctrlrepl_wEna; // @[MCache.scala 86:20]
  wire [31:0] ctrl_io_ctrlrepl_wData; // @[MCache.scala 86:20]
  wire [31:0] ctrl_io_ctrlrepl_wAddr; // @[MCache.scala 86:20]
  wire  ctrl_io_ctrlrepl_wTag; // @[MCache.scala 86:20]
  wire [10:0] ctrl_io_ctrlrepl_addrEven; // @[MCache.scala 86:20]
  wire [10:0] ctrl_io_ctrlrepl_addrOdd; // @[MCache.scala 86:20]
  wire  ctrl_io_ctrlrepl_instrStall; // @[MCache.scala 86:20]
  wire  ctrl_io_replctrl_hit; // @[MCache.scala 86:20]
  wire [31:0] ctrl_io_femcache_addrEven; // @[MCache.scala 86:20]
  wire [31:0] ctrl_io_femcache_addrOdd; // @[MCache.scala 86:20]
  wire  ctrl_io_exmcache_doCallRet; // @[MCache.scala 86:20]
  wire [31:0] ctrl_io_exmcache_callRetBase; // @[MCache.scala 86:20]
  wire [2:0] ctrl_io_ocp_port_M_Cmd; // @[MCache.scala 86:20]
  wire [31:0] ctrl_io_ocp_port_M_Addr; // @[MCache.scala 86:20]
  wire [1:0] ctrl_io_ocp_port_S_Resp; // @[MCache.scala 86:20]
  wire [31:0] ctrl_io_ocp_port_S_Data; // @[MCache.scala 86:20]
  wire  ctrl_io_ocp_port_S_CmdAccept; // @[MCache.scala 86:20]
  wire  ctrl_io_illMem; // @[MCache.scala 86:20]
  wire  ctrl_io_forceHit; // @[MCache.scala 86:20]
  wire  repl_clock; // @[MCache.scala 87:20]
  wire  repl_reset; // @[MCache.scala 87:20]
  wire  repl_io_ena_in; // @[MCache.scala 87:20]
  wire  repl_io_invalidate; // @[MCache.scala 87:20]
  wire  repl_io_hitEna; // @[MCache.scala 87:20]
  wire  repl_io_exmcache_doCallRet; // @[MCache.scala 87:20]
  wire [31:0] repl_io_exmcache_callRetBase; // @[MCache.scala 87:20]
  wire [31:0] repl_io_exmcache_callRetAddr; // @[MCache.scala 87:20]
  wire [31:0] repl_io_mcachefe_instrEven; // @[MCache.scala 87:20]
  wire [31:0] repl_io_mcachefe_instrOdd; // @[MCache.scala 87:20]
  wire [31:0] repl_io_mcachefe_base; // @[MCache.scala 87:20]
  wire [10:0] repl_io_mcachefe_relBase; // @[MCache.scala 87:20]
  wire [11:0] repl_io_mcachefe_relPc; // @[MCache.scala 87:20]
  wire [31:0] repl_io_mcachefe_reloc; // @[MCache.scala 87:20]
  wire [1:0] repl_io_mcachefe_memSel; // @[MCache.scala 87:20]
  wire  repl_io_ctrlrepl_wEna; // @[MCache.scala 87:20]
  wire [31:0] repl_io_ctrlrepl_wData; // @[MCache.scala 87:20]
  wire [31:0] repl_io_ctrlrepl_wAddr; // @[MCache.scala 87:20]
  wire  repl_io_ctrlrepl_wTag; // @[MCache.scala 87:20]
  wire [10:0] repl_io_ctrlrepl_addrEven; // @[MCache.scala 87:20]
  wire [10:0] repl_io_ctrlrepl_addrOdd; // @[MCache.scala 87:20]
  wire  repl_io_ctrlrepl_instrStall; // @[MCache.scala 87:20]
  wire  repl_io_replctrl_hit; // @[MCache.scala 87:20]
  wire  repl_io_memIn_wEven; // @[MCache.scala 87:20]
  wire  repl_io_memIn_wOdd; // @[MCache.scala 87:20]
  wire [31:0] repl_io_memIn_wData; // @[MCache.scala 87:20]
  wire [9:0] repl_io_memIn_wAddr; // @[MCache.scala 87:20]
  wire [9:0] repl_io_memIn_addrEven; // @[MCache.scala 87:20]
  wire [9:0] repl_io_memIn_addrOdd; // @[MCache.scala 87:20]
  wire [31:0] repl_io_memOut_instrEven; // @[MCache.scala 87:20]
  wire [31:0] repl_io_memOut_instrOdd; // @[MCache.scala 87:20]
  wire  mem_clock; // @[MCache.scala 90:19]
  wire  mem_io_memIn_wEven; // @[MCache.scala 90:19]
  wire  mem_io_memIn_wOdd; // @[MCache.scala 90:19]
  wire [31:0] mem_io_memIn_wData; // @[MCache.scala 90:19]
  wire [9:0] mem_io_memIn_wAddr; // @[MCache.scala 90:19]
  wire [9:0] mem_io_memIn_addrEven; // @[MCache.scala 90:19]
  wire [9:0] mem_io_memIn_addrOdd; // @[MCache.scala 90:19]
  wire [31:0] mem_io_memOut_instrEven; // @[MCache.scala 90:19]
  wire [31:0] mem_io_memOut_instrOdd; // @[MCache.scala 90:19]
  MCacheCtrl ctrl ( // @[MCache.scala 86:20]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_fetchEna(ctrl_io_fetchEna),
    .io_ctrlrepl_wEna(ctrl_io_ctrlrepl_wEna),
    .io_ctrlrepl_wData(ctrl_io_ctrlrepl_wData),
    .io_ctrlrepl_wAddr(ctrl_io_ctrlrepl_wAddr),
    .io_ctrlrepl_wTag(ctrl_io_ctrlrepl_wTag),
    .io_ctrlrepl_addrEven(ctrl_io_ctrlrepl_addrEven),
    .io_ctrlrepl_addrOdd(ctrl_io_ctrlrepl_addrOdd),
    .io_ctrlrepl_instrStall(ctrl_io_ctrlrepl_instrStall),
    .io_replctrl_hit(ctrl_io_replctrl_hit),
    .io_femcache_addrEven(ctrl_io_femcache_addrEven),
    .io_femcache_addrOdd(ctrl_io_femcache_addrOdd),
    .io_exmcache_doCallRet(ctrl_io_exmcache_doCallRet),
    .io_exmcache_callRetBase(ctrl_io_exmcache_callRetBase),
    .io_ocp_port_M_Cmd(ctrl_io_ocp_port_M_Cmd),
    .io_ocp_port_M_Addr(ctrl_io_ocp_port_M_Addr),
    .io_ocp_port_S_Resp(ctrl_io_ocp_port_S_Resp),
    .io_ocp_port_S_Data(ctrl_io_ocp_port_S_Data),
    .io_ocp_port_S_CmdAccept(ctrl_io_ocp_port_S_CmdAccept),
    .io_illMem(ctrl_io_illMem),
    .io_forceHit(ctrl_io_forceHit)
  );
  MCacheReplFifo repl ( // @[MCache.scala 87:20]
    .clock(repl_clock),
    .reset(repl_reset),
    .io_ena_in(repl_io_ena_in),
    .io_invalidate(repl_io_invalidate),
    .io_hitEna(repl_io_hitEna),
    .io_exmcache_doCallRet(repl_io_exmcache_doCallRet),
    .io_exmcache_callRetBase(repl_io_exmcache_callRetBase),
    .io_exmcache_callRetAddr(repl_io_exmcache_callRetAddr),
    .io_mcachefe_instrEven(repl_io_mcachefe_instrEven),
    .io_mcachefe_instrOdd(repl_io_mcachefe_instrOdd),
    .io_mcachefe_base(repl_io_mcachefe_base),
    .io_mcachefe_relBase(repl_io_mcachefe_relBase),
    .io_mcachefe_relPc(repl_io_mcachefe_relPc),
    .io_mcachefe_reloc(repl_io_mcachefe_reloc),
    .io_mcachefe_memSel(repl_io_mcachefe_memSel),
    .io_ctrlrepl_wEna(repl_io_ctrlrepl_wEna),
    .io_ctrlrepl_wData(repl_io_ctrlrepl_wData),
    .io_ctrlrepl_wAddr(repl_io_ctrlrepl_wAddr),
    .io_ctrlrepl_wTag(repl_io_ctrlrepl_wTag),
    .io_ctrlrepl_addrEven(repl_io_ctrlrepl_addrEven),
    .io_ctrlrepl_addrOdd(repl_io_ctrlrepl_addrOdd),
    .io_ctrlrepl_instrStall(repl_io_ctrlrepl_instrStall),
    .io_replctrl_hit(repl_io_replctrl_hit),
    .io_memIn_wEven(repl_io_memIn_wEven),
    .io_memIn_wOdd(repl_io_memIn_wOdd),
    .io_memIn_wData(repl_io_memIn_wData),
    .io_memIn_wAddr(repl_io_memIn_wAddr),
    .io_memIn_addrEven(repl_io_memIn_addrEven),
    .io_memIn_addrOdd(repl_io_memIn_addrOdd),
    .io_memOut_instrEven(repl_io_memOut_instrEven),
    .io_memOut_instrOdd(repl_io_memOut_instrOdd)
  );
  MCacheMem mem ( // @[MCache.scala 90:19]
    .clock(mem_clock),
    .io_memIn_wEven(mem_io_memIn_wEven),
    .io_memIn_wOdd(mem_io_memIn_wOdd),
    .io_memIn_wData(mem_io_memIn_wData),
    .io_memIn_wAddr(mem_io_memIn_wAddr),
    .io_memIn_addrEven(mem_io_memIn_addrEven),
    .io_memIn_addrOdd(mem_io_memIn_addrOdd),
    .io_memOut_instrEven(mem_io_memOut_instrEven),
    .io_memOut_instrOdd(mem_io_memOut_instrOdd)
  );
  assign io_ena_out = ctrl_io_fetchEna & (repl_io_hitEna | ctrl_io_forceHit); // @[MCache.scala 108:34]
  assign io_icachefe_instrEven = repl_io_mcachefe_instrEven; // @[MCache.scala 98:15]
  assign io_icachefe_instrOdd = repl_io_mcachefe_instrOdd; // @[MCache.scala 98:15]
  assign io_icachefe_base = repl_io_mcachefe_base; // @[MCache.scala 98:15]
  assign io_icachefe_relBase = repl_io_mcachefe_relBase; // @[MCache.scala 98:15]
  assign io_icachefe_relPc = repl_io_mcachefe_relPc; // @[MCache.scala 98:15]
  assign io_icachefe_reloc = repl_io_mcachefe_reloc; // @[MCache.scala 98:15]
  assign io_icachefe_memSel = repl_io_mcachefe_memSel; // @[MCache.scala 98:15]
  assign io_ocp_port_M_Cmd = ctrl_io_ocp_port_M_Cmd; // @[MCache.scala 95:15]
  assign io_ocp_port_M_Addr = ctrl_io_ocp_port_M_Addr; // @[MCache.scala 95:15]
  assign io_illMem = ctrl_io_illMem; // @[MCache.scala 110:13]
  assign ctrl_clock = clock;
  assign ctrl_reset = reset;
  assign ctrl_io_replctrl_hit = repl_io_replctrl_hit; // @[MCache.scala 99:20]
  assign ctrl_io_femcache_addrEven = io_feicache_addrEven; // @[MCache.scala 93:20]
  assign ctrl_io_femcache_addrOdd = io_feicache_addrOdd; // @[MCache.scala 93:20]
  assign ctrl_io_exmcache_doCallRet = io_exicache_doCallRet; // @[MCache.scala 94:20]
  assign ctrl_io_exmcache_callRetBase = io_exicache_callRetBase; // @[MCache.scala 94:20]
  assign ctrl_io_ocp_port_S_Resp = io_ocp_port_S_Resp; // @[MCache.scala 95:15]
  assign ctrl_io_ocp_port_S_Data = io_ocp_port_S_Data; // @[MCache.scala 95:15]
  assign ctrl_io_ocp_port_S_CmdAccept = io_ocp_port_S_CmdAccept; // @[MCache.scala 95:15]
  assign repl_clock = clock;
  assign repl_reset = reset;
  assign repl_io_ena_in = io_ena_in; // @[MCache.scala 106:18]
  assign repl_io_invalidate = io_invalidate | ctrl_io_illMem; // @[MCache.scala 112:39]
  assign repl_io_exmcache_doCallRet = io_exicache_doCallRet; // @[MCache.scala 97:20]
  assign repl_io_exmcache_callRetBase = io_exicache_callRetBase; // @[MCache.scala 97:20]
  assign repl_io_exmcache_callRetAddr = io_exicache_callRetAddr; // @[MCache.scala 97:20]
  assign repl_io_ctrlrepl_wEna = ctrl_io_ctrlrepl_wEna; // @[MCache.scala 92:20]
  assign repl_io_ctrlrepl_wData = ctrl_io_ctrlrepl_wData; // @[MCache.scala 92:20]
  assign repl_io_ctrlrepl_wAddr = ctrl_io_ctrlrepl_wAddr; // @[MCache.scala 92:20]
  assign repl_io_ctrlrepl_wTag = ctrl_io_ctrlrepl_wTag; // @[MCache.scala 92:20]
  assign repl_io_ctrlrepl_addrEven = ctrl_io_ctrlrepl_addrEven; // @[MCache.scala 92:20]
  assign repl_io_ctrlrepl_addrOdd = ctrl_io_ctrlrepl_addrOdd; // @[MCache.scala 92:20]
  assign repl_io_ctrlrepl_instrStall = ctrl_io_ctrlrepl_instrStall; // @[MCache.scala 92:20]
  assign repl_io_memOut_instrEven = mem_io_memOut_instrEven; // @[MCache.scala 103:18]
  assign repl_io_memOut_instrOdd = mem_io_memOut_instrOdd; // @[MCache.scala 103:18]
  assign mem_clock = clock;
  assign mem_io_memIn_wEven = repl_io_memIn_wEven; // @[MCache.scala 102:16]
  assign mem_io_memIn_wOdd = repl_io_memIn_wOdd; // @[MCache.scala 102:16]
  assign mem_io_memIn_wData = repl_io_memIn_wData; // @[MCache.scala 102:16]
  assign mem_io_memIn_wAddr = repl_io_memIn_wAddr; // @[MCache.scala 102:16]
  assign mem_io_memIn_addrEven = repl_io_memIn_addrEven; // @[MCache.scala 102:16]
  assign mem_io_memIn_addrOdd = repl_io_memIn_addrOdd; // @[MCache.scala 102:16]
endmodule
module MemBlock_2(
  input         clock,
  input  [6:0]  io_rdAddr,
  output [31:0] io_rdData,
  input  [6:0]  io_wrAddr,
  input         io_wrEna,
  input  [31:0] io_wrData
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:127];
  wire [31:0] mem_MPORT_1_data;
  wire [6:0] mem_MPORT_1_addr;
  wire [31:0] mem_MPORT_data;
  wire [6:0] mem_MPORT_addr;
  wire  mem_MPORT_mask;
  wire  mem_MPORT_en;
  reg [6:0] rdAddrReg; // @[MemBlock.scala 59:22]
  assign mem_MPORT_1_addr = rdAddrReg;
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr];
  assign mem_MPORT_data = io_wrData;
  assign mem_MPORT_addr = io_wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEna;
  assign io_rdData = mem_MPORT_1_data; // @[MemBlock.scala 60:13]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data;
    end
    rdAddrReg <= io_rdAddr; // @[MemBlock.scala 59:22]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rdAddrReg = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Fetch(
  input         clock,
  input         reset,
  input         io_ena,
  output [31:0] io_fedec_instr_a,
  output [31:0] io_fedec_instr_b,
  output [29:0] io_fedec_pc,
  output [29:0] io_fedec_base,
  output [31:0] io_fedec_reloc,
  output [29:0] io_fedec_relPc,
  output [29:0] io_feex_pc,
  input         io_exfe_doBranch,
  input  [29:0] io_exfe_branchPc,
  input         io_memfe_doCallRet,
  input         io_memfe_store,
  input  [31:0] io_memfe_addr,
  input  [31:0] io_memfe_data,
  output [31:0] io_feicache_addrEven,
  output [31:0] io_feicache_addrOdd,
  input  [31:0] io_icachefe_instrEven,
  input  [31:0] io_icachefe_instrOdd,
  input  [31:0] io_icachefe_base,
  input  [10:0] io_icachefe_relBase,
  input  [11:0] io_icachefe_relPc,
  input  [31:0] io_icachefe_reloc,
  input  [1:0]  io_icachefe_memSel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  MemBlock_clock; // @[MemBlock.scala 15:11]
  wire [6:0] MemBlock_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [31:0] MemBlock_io_rdData; // @[MemBlock.scala 15:11]
  wire [6:0] MemBlock_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_io_wrEna; // @[MemBlock.scala 15:11]
  wire [31:0] MemBlock_io_wrData; // @[MemBlock.scala 15:11]
  wire  MemBlock_1_clock; // @[MemBlock.scala 15:11]
  wire [6:0] MemBlock_1_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [31:0] MemBlock_1_io_rdData; // @[MemBlock.scala 15:11]
  wire [6:0] MemBlock_1_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_1_io_wrEna; // @[MemBlock.scala 15:11]
  wire [31:0] MemBlock_1_io_wrData; // @[MemBlock.scala 15:11]
  reg [29:0] pcReg; // @[Fetch.scala 21:22]
  reg [29:0] addrEvenReg; // @[Fetch.scala 25:24]
  reg [29:0] addrOddReg; // @[Fetch.scala 26:23]
  wire  _T_2 = io_memfe_store & io_memfe_addr[31:16] == 16'h1; // @[Fetch.scala 48:36]
  reg  selSpm; // @[Fetch.scala 65:23]
  wire  _T_14 = ~pcReg[0]; // @[Fetch.scala 57:34]
  wire [31:0] instr_a_ispm = ~pcReg[0] ? MemBlock_io_rdData : MemBlock_1_io_rdData; // @[Fetch.scala 57:24]
  reg  selCache; // @[Fetch.scala 66:25]
  wire [31:0] instr_a_cache = _T_14 ? io_icachefe_instrEven : io_icachefe_instrOdd; // @[Fetch.scala 106:26]
  reg [31:0] data_even; // @[Fetch.scala 100:26]
  reg [31:0] data_odd; // @[Fetch.scala 101:25]
  wire [31:0] instr_a_rom = _T_14 ? data_even : data_odd; // @[Fetch.scala 102:24]
  wire [31:0] _T_31 = selCache ? instr_a_cache : instr_a_rom; // @[Fetch.scala 111:24]
  wire [31:0] instr_a = selSpm ? instr_a_ispm : _T_31; // @[Fetch.scala 110:20]
  wire  b_valid = instr_a[31]; // @[Fetch.scala 115:24]
  wire [29:0] _T_35 = pcReg + 30'h2; // @[Fetch.scala 117:36]
  wire [29:0] _T_37 = pcReg + 30'h1; // @[Fetch.scala 117:53]
  wire [29:0] pc_cont = b_valid ? _T_35 : _T_37; // @[Fetch.scala 117:20]
  wire [29:0] _T_38 = io_exfe_doBranch ? io_exfe_branchPc : pc_cont; // @[Fetch.scala 120:16]
  wire [29:0] pc_next = io_memfe_doCallRet ? {{18'd0}, io_icachefe_relPc} : _T_38; // @[Fetch.scala 119:8]
  wire [11:0] _T_44 = io_icachefe_relPc + 12'h2; // @[Fetch.scala 125:54]
  wire [29:0] _T_46 = io_exfe_branchPc + 30'h2; // @[Fetch.scala 126:48]
  wire [29:0] _T_40 = pcReg + 30'h4; // @[Fetch.scala 123:37]
  wire [29:0] _T_42 = pcReg + 30'h3; // @[Fetch.scala 123:54]
  wire [29:0] pc_cont2 = b_valid ? _T_40 : _T_42; // @[Fetch.scala 123:21]
  wire [29:0] _T_47 = io_exfe_doBranch ? _T_46 : pc_cont2; // @[Fetch.scala 126:12]
  wire [29:0] pc_next2 = io_memfe_doCallRet ? {{18'd0}, _T_44} : _T_47; // @[Fetch.scala 125:8]
  wire [29:0] pc_inc = pc_next[0] ? pc_next2 : pc_next; // @[Fetch.scala 129:19]
  wire [28:0] hi = pc_inc[29:1]; // @[Fetch.scala 133:29]
  wire [29:0] _T_52 = {hi,1'h0}; // @[Cat.scala 30:58]
  wire [29:0] addrEven = io_ena & ~reset ? _T_52 : addrEvenReg; // @[Fetch.scala 132:26 Fetch.scala 133:14 Fetch.scala 130:12]
  wire [28:0] hi_1 = pc_next[29:1]; // @[Fetch.scala 134:29]
  wire [29:0] _T_53 = {hi_1,1'h1}; // @[Cat.scala 30:58]
  wire [29:0] addrOdd = io_ena & ~reset ? _T_53 : addrOddReg; // @[Fetch.scala 132:26 Fetch.scala 134:13 Fetch.scala 131:11]
  wire [31:0] instr_b_ispm = _T_14 ? MemBlock_1_io_rdData : MemBlock_io_rdData; // @[Fetch.scala 58:24]
  reg [31:0] baseReg; // @[Fetch.scala 79:24]
  reg [10:0] relBaseReg; // @[Fetch.scala 80:27]
  reg [31:0] relocReg; // @[Fetch.scala 81:25]
  wire [10:0] _GEN_2 = io_memfe_doCallRet ? io_icachefe_relBase : relBaseReg; // @[Fetch.scala 91:31 Fetch.scala 92:19 Fetch.scala 85:15]
  wire [31:0] _GEN_3 = io_memfe_doCallRet ? io_icachefe_reloc : relocReg; // @[Fetch.scala 91:31 Fetch.scala 93:17 Fetch.scala 87:13]
  wire [31:0] _GEN_8 = 9'h1 == addrEven[9:1] ? 32'h20700 : 32'h54; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_9 = 9'h2 == addrEven[9:1] ? 32'h20800 : _GEN_8; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_10 = 9'h3 == addrEven[9:1] ? 32'h2402025 : _GEN_9; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_11 = 9'h4 == addrEven[9:1] ? 32'h87c20000 : _GEN_10; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_12 = 9'h5 == addrEven[9:1] ? 32'h2821085 : _GEN_11; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_13 = 9'h6 == addrEven[9:1] ? 32'h2021062 : _GEN_12; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_14 = 9'h7 == addrEven[9:1] ? 32'hf0010000 : _GEN_13; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_15 = 9'h8 == addrEven[9:1] ? 32'h80000000 : _GEN_14; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_16 = 9'h9 == addrEven[9:1] ? 32'h400000 : _GEN_15; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_17 = 9'ha == addrEven[9:1] ? 32'h4000017 : _GEN_16; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_18 = 9'hb == addrEven[9:1] ? 32'h4ac : _GEN_17; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_19 = 9'hc == addrEven[9:1] ? 32'h2520038 : _GEN_18; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_20 = 9'hd == addrEven[9:1] ? 32'h2c5fd08 : _GEN_19; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_21 = 9'he == addrEven[9:1] ? 32'h2c5f481 : _GEN_20; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_22 = 9'hf == addrEven[9:1] ? 32'h2c5f480 : _GEN_21; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_23 = 9'h10 == addrEven[9:1] ? 32'h2c5fb04 : _GEN_22; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_24 = 9'h11 == addrEven[9:1] ? 32'h2c5fc06 : _GEN_23; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_25 = 9'h12 == addrEven[9:1] ? 32'h87c20000 : _GEN_24; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_26 = 9'h13 == addrEven[9:1] ? 32'h2821083 : _GEN_25; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_27 = 9'h14 == addrEven[9:1] ? 32'h2022081 : _GEN_26; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_28 = 9'h15 == addrEven[9:1] ? 32'hf0020000 : _GEN_27; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_29 = 9'h16 == addrEven[9:1] ? 32'h400000 : _GEN_28; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_30 = 9'h17 == addrEven[9:1] ? 32'h2022062 : _GEN_29; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_31 = 9'h18 == addrEven[9:1] ? 32'h2c60005 : _GEN_30; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_32 = 9'h19 == addrEven[9:1] ? 32'h87c20000 : _GEN_31; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_33 = 9'h1a == addrEven[9:1] ? 32'h2821080 : _GEN_32; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_34 = 9'h1b == addrEven[9:1] ? 32'h2021031 : _GEN_33; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_35 = 9'h1c == addrEven[9:1] ? 32'h87c20000 : _GEN_34; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_36 = 9'h1d == addrEven[9:1] ? 32'h2841080 : _GEN_35; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_37 = 9'h1e == addrEven[9:1] ? 32'hc42004 : _GEN_36; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_38 = 9'h1f == addrEven[9:1] ? 32'h2841080 : _GEN_37; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_39 = 9'h20 == addrEven[9:1] ? 32'hc42004 : _GEN_38; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_40 = 9'h21 == addrEven[9:1] ? 32'h2841080 : _GEN_39; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_41 = 9'h22 == addrEven[9:1] ? 32'hc42004 : _GEN_40; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_42 = 9'h23 == addrEven[9:1] ? 32'h2821080 : _GEN_41; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_43 = 9'h24 == addrEven[9:1] ? 32'hc21004 : _GEN_42; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_44 = 9'h25 == addrEven[9:1] ? 32'h40001 : _GEN_43; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_45 = 9'h26 == addrEven[9:1] ? 32'hf0000000 : _GEN_44; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_46 = 9'h27 == addrEven[9:1] ? 32'h400000 : _GEN_45; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_47 = 9'h28 == addrEven[9:1] ? 32'h2c61109 : _GEN_46; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_48 = 9'h29 == addrEven[9:1] ? 32'h400000 : _GEN_47; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_49 = 9'h2a == addrEven[9:1] ? 32'hcbffff7 : _GEN_48; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_50 = 9'h2b == addrEven[9:1] ? 32'h400000 : _GEN_49; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_51 = 9'h2c == addrEven[9:1] ? 32'hcbffffd : _GEN_50; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_52 = 9'h2d == addrEven[9:1] ? 32'h87c40000 : _GEN_51; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_53 = 9'h2e == addrEven[9:1] ? 32'h2842082 : _GEN_52; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_54 = 9'h2f == addrEven[9:1] ? 32'h2022060 : _GEN_53; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_55 = 9'h30 == addrEven[9:1] ? 32'h20010 : _GEN_54; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_56 = 9'h31 == addrEven[9:1] ? 32'hc22004 : _GEN_55; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_57 = 9'h32 == addrEven[9:1] ? 32'h460001 : _GEN_56; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_58 = 9'h33 == addrEven[9:1] ? 32'h2c61007 : _GEN_57; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_59 = 9'h34 == addrEven[9:1] ? 32'h20010 : _GEN_58; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_60 = 9'h35 == addrEven[9:1] ? 32'hf0000000 : _GEN_59; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_61 = 9'h36 == addrEven[9:1] ? 32'h42001 : _GEN_60; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_62 = 9'h37 == addrEven[9:1] ? 32'hcbffff4 : _GEN_61; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_63 = 9'h38 == addrEven[9:1] ? 32'h2021031 : _GEN_62; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_64 = 9'h39 == addrEven[9:1] ? 32'h40001 : _GEN_63; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_65 = 9'h3a == addrEven[9:1] ? 32'h4000143 : _GEN_64; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_66 = 9'h3b == addrEven[9:1] ? 32'h87c20000 : _GEN_65; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_67 = 9'h3c == addrEven[9:1] ? 32'h282108c : _GEN_66; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_68 = 9'h3d == addrEven[9:1] ? 32'h2021264 : _GEN_67; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_69 = 9'h3e == addrEven[9:1] ? 32'hc80000d : _GEN_68; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_70 = 9'h3f == addrEven[9:1] ? 32'h10000 : _GEN_69; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_71 = 9'h40 == addrEven[9:1] ? 32'h400000 : _GEN_70; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_72 = 9'h41 == addrEven[9:1] ? 32'h87c40000 : _GEN_71; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_73 = 9'h42 == addrEven[9:1] ? 32'h284208c : _GEN_72; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_74 = 9'h43 == addrEven[9:1] ? 32'h1042002 : _GEN_73; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_75 = 9'h44 == addrEven[9:1] ? 32'hcbffff5 : _GEN_74; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_76 = 9'h45 == addrEven[9:1] ? 32'hf0000000 : _GEN_75; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_77 = 9'h46 == addrEven[9:1] ? 32'h400000 : _GEN_76; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_78 = 9'h47 == addrEven[9:1] ? 32'h4c800008 : _GEN_77; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_79 = 9'h48 == addrEven[9:1] ? 32'hf0000000 : _GEN_78; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_80 = 9'h49 == addrEven[9:1] ? 32'h40002 : _GEN_79; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_81 = 9'h4a == addrEven[9:1] ? 32'hc21004 : _GEN_80; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_82 = 9'h4b == addrEven[9:1] ? 32'h20002 : _GEN_81; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_83 = 9'h4c == addrEven[9:1] ? 32'h87c40000 : _GEN_82; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_84 = 9'h4d == addrEven[9:1] ? 32'h2842082 : _GEN_83; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_85 = 9'h4e == addrEven[9:1] ? 32'h2022164 : _GEN_84; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_86 = 9'h4f == addrEven[9:1] ? 32'hc41004 : _GEN_85; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_87 = 9'h50 == addrEven[9:1] ? 32'h400000 : _GEN_86; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_88 = 9'h51 == addrEven[9:1] ? 32'hcbffffc : _GEN_87; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_89 = 9'h52 == addrEven[9:1] ? 32'hf0000000 : _GEN_88; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_90 = 9'h53 == addrEven[9:1] ? 32'h21001 : _GEN_89; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_91 = 9'h54 == addrEven[9:1] ? 32'hcbffff6 : _GEN_90; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_92 = 9'h55 == addrEven[9:1] ? 32'h200ff : _GEN_91; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_93 = 9'h56 == addrEven[9:1] ? 32'hc800023 : _GEN_92; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_94 = 9'h57 == addrEven[9:1] ? 32'hf0010000 : _GEN_93; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_95 = 9'h58 == addrEven[9:1] ? 32'h440001 : _GEN_94; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_96 = 9'h59 == addrEven[9:1] ? 32'hcfc40000 : _GEN_95; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_97 = 9'h5a == addrEven[9:1] ? 32'hcfc20000 : _GEN_96; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_98 = 9'h5b == addrEven[9:1] ? 32'h4ac22085 : _GEN_97; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_99 = 9'h5c == addrEven[9:1] ? 32'h400000 : _GEN_98; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_100 = 9'h5d == addrEven[9:1] ? 32'h400000 : _GEN_99; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_101 = 9'h5e == addrEven[9:1] ? 32'h87c40000 : _GEN_100; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_102 = 9'h5f == addrEven[9:1] ? 32'h2842085 : _GEN_101; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_103 = 9'h60 == addrEven[9:1] ? 32'h2022062 : _GEN_102; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_104 = 9'h61 == addrEven[9:1] ? 32'hf0010000 : _GEN_103; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_105 = 9'h62 == addrEven[9:1] ? 32'h80000000 : _GEN_104; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_106 = 9'h63 == addrEven[9:1] ? 32'h400000 : _GEN_105; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_107 = 9'h64 == addrEven[9:1] ? 32'h87c40000 : _GEN_106; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_108 = 9'h65 == addrEven[9:1] ? 32'h2842080 : _GEN_107; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_109 = 9'h66 == addrEven[9:1] ? 32'hc42004 : _GEN_108; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_110 = 9'h67 == addrEven[9:1] ? 32'h1c210ff : _GEN_109; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_111 = 9'h68 == addrEven[9:1] ? 32'hf0000000 : _GEN_110; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_112 = 9'h69 == addrEven[9:1] ? 32'h400000 : _GEN_111; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_113 = 9'h6a == addrEven[9:1] ? 32'h4c800012 : _GEN_112; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_114 = 9'h6b == addrEven[9:1] ? 32'h87c20000 : _GEN_113; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_115 = 9'h6c == addrEven[9:1] ? 32'h2821080 : _GEN_114; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_116 = 9'h6d == addrEven[9:1] ? 32'hc21004 : _GEN_115; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_117 = 9'h6e == addrEven[9:1] ? 32'h2820185 : _GEN_116; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_118 = 9'h6f == addrEven[9:1] ? 32'h2021261 : _GEN_117; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_119 = 9'h70 == addrEven[9:1] ? 32'h87c20000 : _GEN_118; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_120 = 9'h71 == addrEven[9:1] ? 32'h2821080 : _GEN_119; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_121 = 9'h72 == addrEven[9:1] ? 32'hc21004 : _GEN_120; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_122 = 9'h73 == addrEven[9:1] ? 32'h87c60000 : _GEN_121; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_123 = 9'h74 == addrEven[9:1] ? 32'h2863082 : _GEN_122; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_124 = 9'h75 == addrEven[9:1] ? 32'h2023164 : _GEN_123; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_125 = 9'h76 == addrEven[9:1] ? 32'hc62004 : _GEN_124; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_126 = 9'h77 == addrEven[9:1] ? 32'h400000 : _GEN_125; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_127 = 9'h78 == addrEven[9:1] ? 32'hc800006 : _GEN_126; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_128 = 9'h79 == addrEven[9:1] ? 32'h2863189 : _GEN_127; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_129 = 9'h7a == addrEven[9:1] ? 32'h2023261 : _GEN_128; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_130 = 9'h7b == addrEven[9:1] ? 32'h87c60000 : _GEN_129; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_131 = 9'h7c == addrEven[9:1] ? 32'h2863082 : _GEN_130; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_132 = 9'h7d == addrEven[9:1] ? 32'h20221b4 : _GEN_131; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_133 = 9'h7e == addrEven[9:1] ? 32'h87c40000 : _GEN_132; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_134 = 9'h7f == addrEven[9:1] ? 32'h2842080 : _GEN_133; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_135 = 9'h80 == addrEven[9:1] ? 32'h2022036 : _GEN_134; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_136 = 9'h81 == addrEven[9:1] ? 32'h87c40000 : _GEN_135; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_137 = 9'h82 == addrEven[9:1] ? 32'h2c22001 : _GEN_136; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_138 = 9'h83 == addrEven[9:1] ? 32'hf0080000 : _GEN_137; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_139 = 9'h84 == addrEven[9:1] ? 32'h400000 : _GEN_138; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_140 = 9'h85 == addrEven[9:1] ? 32'h4cbffffb : _GEN_139; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_141 = 9'h86 == addrEven[9:1] ? 32'h87c60000 : _GEN_140; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_142 = 9'h87 == addrEven[9:1] ? 32'h2c23101 : _GEN_141; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_143 = 9'h88 == addrEven[9:1] ? 32'hf0080000 : _GEN_142; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_144 = 9'h89 == addrEven[9:1] ? 32'h400000 : _GEN_143; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_145 = 9'h8a == addrEven[9:1] ? 32'h4cbffffb : _GEN_144; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_146 = 9'h8b == addrEven[9:1] ? 32'hf0080000 : _GEN_145; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_147 = 9'h8c == addrEven[9:1] ? 32'h20004 : _GEN_146; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_148 = 9'h8d == addrEven[9:1] ? 32'h87c40000 : _GEN_147; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_149 = 9'h8e == addrEven[9:1] ? 32'h2842082 : _GEN_148; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_150 = 9'h8f == addrEven[9:1] ? 32'h2022164 : _GEN_149; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_151 = 9'h90 == addrEven[9:1] ? 32'hc41004 : _GEN_150; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_152 = 9'h91 == addrEven[9:1] ? 32'h400000 : _GEN_151; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_153 = 9'h92 == addrEven[9:1] ? 32'hcbffffc : _GEN_152; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_154 = 9'h93 == addrEven[9:1] ? 32'hf0000000 : _GEN_153; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_155 = 9'h94 == addrEven[9:1] ? 32'h21001 : _GEN_154; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_156 = 9'h95 == addrEven[9:1] ? 32'hcbffff6 : _GEN_155; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_157 = 9'h96 == addrEven[9:1] ? 32'hf0010000 : _GEN_156; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_158 = 9'h97 == addrEven[9:1] ? 32'h4400001 : _GEN_157; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_159 = 9'h98 == addrEven[9:1] ? 32'h20002 : _GEN_158; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_160 = 9'h99 == addrEven[9:1] ? 32'h2adf104 : _GEN_159; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_161 = 9'h9a == addrEven[9:1] ? 32'h2b1f106 : _GEN_160; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_162 = 9'h9b == addrEven[9:1] ? 32'h2b5f108 : _GEN_161; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_163 = 9'h9c == addrEven[9:1] ? 32'h2abf103 : _GEN_162; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_164 = 9'h9d == addrEven[9:1] ? 32'h293f101 : _GEN_163; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_165 = 9'h9e == addrEven[9:1] ? 32'h2409027 : _GEN_164; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_166 = 9'h9f == addrEven[9:1] ? 32'h6400000 : _GEN_165; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_167 = 9'ha0 == addrEven[9:1] ? 32'h2409020 : _GEN_166; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_168 = 9'ha1 == addrEven[9:1] ? 32'h340 : _GEN_167; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_169 = 9'ha2 == addrEven[9:1] ? 32'h2520038 : _GEN_168; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_170 = 9'ha3 == addrEven[9:1] ? 32'h87c20000 : _GEN_169; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_171 = 9'ha4 == addrEven[9:1] ? 32'h2c41000 : _GEN_170; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_172 = 9'ha5 == addrEven[9:1] ? 32'h2520037 : _GEN_171; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_173 = 9'ha6 == addrEven[9:1] ? 32'h2520030 : _GEN_172; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_174 = 9'ha7 == addrEven[9:1] ? 32'h2c5fa88 : _GEN_173; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_175 = 9'ha8 == addrEven[9:1] ? 32'h2c5fb8a : _GEN_174; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_176 = 9'ha9 == addrEven[9:1] ? 32'h2c5fc8c : _GEN_175; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_177 = 9'haa == addrEven[9:1] ? 32'h2c5fd8e : _GEN_176; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_178 = 9'hab == addrEven[9:1] ? 32'h87c21000 : _GEN_177; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_179 = 9'hac == addrEven[9:1] ? 32'h40020 : _GEN_178; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_180 = 9'had == addrEven[9:1] ? 32'h87c40000 : _GEN_179; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_181 = 9'hae == addrEven[9:1] ? 32'h2822100 : _GEN_180; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_182 = 9'haf == addrEven[9:1] ? 32'h21001 : _GEN_181; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_183 = 9'hb0 == addrEven[9:1] ? 32'h403be : _GEN_182; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_184 = 9'hb1 == addrEven[9:1] ? 32'hcbffff4 : _GEN_183; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_185 = 9'hb2 == addrEven[9:1] ? 32'h20404 : _GEN_184; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_186 = 9'hb3 == addrEven[9:1] ? 32'h460001 : _GEN_185; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_187 = 9'hb4 == addrEven[9:1] ? 32'h360000 : _GEN_186; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_188 = 9'hb5 == addrEven[9:1] ? 32'h2a0000 : _GEN_187; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_189 = 9'hb6 == addrEven[9:1] ? 32'h300000 : _GEN_188; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_190 = 9'hb7 == addrEven[9:1] ? 32'h2c5f000 : _GEN_189; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_191 = 9'hb8 == addrEven[9:1] ? 32'h87c20000 : _GEN_190; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_192 = 9'hb9 == addrEven[9:1] ? 32'h2c41000 : _GEN_191; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_193 = 9'hba == addrEven[9:1] ? 32'h2c5f084 : _GEN_192; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_194 = 9'hbb == addrEven[9:1] ? 32'h20000 : _GEN_193; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_195 = 9'hbc == addrEven[9:1] ? 32'h322000 : _GEN_194; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_196 = 9'hbd == addrEven[9:1] ? 32'h4400214 : _GEN_195; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_197 = 9'hbe == addrEven[9:1] ? 32'hf0090000 : _GEN_196; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_198 = 9'hbf == addrEven[9:1] ? 32'h2c4000 : _GEN_197; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_199 = 9'hc0 == addrEven[9:1] ? 32'h203c060 : _GEN_198; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_200 = 9'hc1 == addrEven[9:1] ? 32'h80000 : _GEN_199; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_201 = 9'hc2 == addrEven[9:1] ? 32'h40003 : _GEN_200; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_202 = 9'hc3 == addrEven[9:1] ? 32'hc800005 : _GEN_201; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_203 = 9'hc4 == addrEven[9:1] ? 32'h4c0005d : _GEN_202; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_204 = 9'hc5 == addrEven[9:1] ? 32'h59000 : _GEN_203; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_205 = 9'hc6 == addrEven[9:1] ? 32'h2022b35 : _GEN_204; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_206 = 9'hc7 == addrEven[9:1] ? 32'h2081c82 : _GEN_205; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_207 = 9'hc8 == addrEven[9:1] ? 32'h1044001 : _GEN_206; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_208 = 9'hc9 == addrEven[9:1] ? 32'h87c42002 : _GEN_207; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_209 = 9'hca == addrEven[9:1] ? 32'h202104a : _GEN_208; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_210 = 9'hcb == addrEven[9:1] ? 32'h82000 : _GEN_209; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_211 = 9'hcc == addrEven[9:1] ? 32'h2023031 : _GEN_210; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_212 = 9'hcd == addrEven[9:1] ? 32'hc75003 : _GEN_211; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_213 = 9'hce == addrEven[9:1] ? 32'h1c63018 : _GEN_212; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_214 = 9'hcf == addrEven[9:1] ? 32'h2021183 : _GEN_213; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_215 = 9'hd0 == addrEven[9:1] ? 32'h20004 : _GEN_214; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_216 = 9'hd1 == addrEven[9:1] ? 32'hcc00013 : _GEN_215; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_217 = 9'hd2 == addrEven[9:1] ? 32'h75001 : _GEN_216; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_218 = 9'hd3 == addrEven[9:1] ? 32'hc800013 : _GEN_217; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_219 = 9'hd4 == addrEven[9:1] ? 32'h2021db4 : _GEN_218; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_220 = 9'hd5 == addrEven[9:1] ? 32'h87c3b00d : _GEN_219; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_221 = 9'hd6 == addrEven[9:1] ? 32'h2861100 : _GEN_220; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_222 = 9'hd7 == addrEven[9:1] ? 32'h6003005 : _GEN_221; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_223 = 9'hd8 == addrEven[9:1] ? 32'h400000 : _GEN_222; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_224 = 9'hd9 == addrEven[9:1] ? 32'h4c00033 : _GEN_223; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_225 = 9'hda == addrEven[9:1] ? 32'h77000 : _GEN_224; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_226 = 9'hdb == addrEven[9:1] ? 32'h87c21007 : _GEN_225; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_227 = 9'hdc == addrEven[9:1] ? 32'h2c61280 : _GEN_226; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_228 = 9'hdd == addrEven[9:1] ? 32'h283f101 : _GEN_227; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_229 = 9'hde == addrEven[9:1] ? 32'h85000 : _GEN_228; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_230 = 9'hdf == addrEven[9:1] ? 32'h305000 : _GEN_229; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_231 = 9'he0 == addrEven[9:1] ? 32'h345000 : _GEN_230; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_232 = 9'he1 == addrEven[9:1] ? 32'h400000 : _GEN_231; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_233 = 9'he2 == addrEven[9:1] ? 32'h60000 : _GEN_232; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_234 = 9'he3 == addrEven[9:1] ? 32'h205b2e0 : _GEN_233; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_235 = 9'he4 == addrEven[9:1] ? 32'h4c800015 : _GEN_234; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_236 = 9'he5 == addrEven[9:1] ? 32'h87c63007 : _GEN_235; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_237 = 9'he6 == addrEven[9:1] ? 32'h203a1b5 : _GEN_236; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_238 = 9'he7 == addrEven[9:1] ? 32'h400000 : _GEN_237; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_239 = 9'he8 == addrEven[9:1] ? 32'h2098180 : _GEN_238; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_240 = 9'he9 == addrEven[9:1] ? 32'h2023d34 : _GEN_239; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_241 = 9'hea == addrEven[9:1] ? 32'h87c84007 : _GEN_240; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_242 = 9'heb == addrEven[9:1] ? 32'h2c64000 : _GEN_241; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_243 = 9'hec == addrEven[9:1] ? 32'h2a0000 : _GEN_242; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_244 = 9'hed == addrEven[9:1] ? 32'h4c00005 : _GEN_243; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_245 = 9'hee == addrEven[9:1] ? 32'h2c5f180 : _GEN_244; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_246 = 9'hef == addrEven[9:1] ? 32'h2a3000 : _GEN_245; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_247 = 9'hf0 == addrEven[9:1] ? 32'h2023060 : _GEN_246; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_248 = 9'hf1 == addrEven[9:1] ? 32'h2c5f283 : _GEN_247; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_249 = 9'hf2 == addrEven[9:1] ? 32'h77000 : _GEN_248; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_250 = 9'hf3 == addrEven[9:1] ? 32'h20360b1 : _GEN_249; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_251 = 9'hf4 == addrEven[9:1] ? 32'h96001 : _GEN_250; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_252 = 9'hf5 == addrEven[9:1] ? 32'h87c20000 : _GEN_251; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_253 = 9'hf6 == addrEven[9:1] ? 32'h2821080 : _GEN_252; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_254 = 9'hf7 == addrEven[9:1] ? 32'h2021036 : _GEN_253; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_255 = 9'hf8 == addrEven[9:1] ? 32'h202200b : _GEN_254; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_256 = 9'hf9 == addrEven[9:1] ? 32'h87ca0000 : _GEN_255; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_257 = 9'hfa == addrEven[9:1] ? 32'h20230b1 : _GEN_256; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_258 = 9'hfb == addrEven[9:1] ? 32'h2c25101 : _GEN_257; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_259 = 9'hfc == addrEven[9:1] ? 32'h283f100 : _GEN_258; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_260 = 9'hfd == addrEven[9:1] ? 32'h400000 : _GEN_259; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_261 = 9'hfe == addrEven[9:1] ? 32'hcffff7b : _GEN_260; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_262 = 9'hff == addrEven[9:1] ? 32'h43000 : _GEN_261; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_263 = 9'h100 == addrEven[9:1] ? 32'h400000 : _GEN_262; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_264 = 9'h101 == addrEven[9:1] ? 32'h2aff10a : _GEN_263; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_265 = 9'h102 == addrEven[9:1] ? 32'h2b3f10c : _GEN_264; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_266 = 9'h103 == addrEven[9:1] ? 32'h2b7f10e : _GEN_265; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_267 = 9'h104 == addrEven[9:1] ? 32'h293f107 : _GEN_266; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_268 = 9'h105 == addrEven[9:1] ? 32'h2409028 : _GEN_267; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_269 = 9'h106 == addrEven[9:1] ? 32'h400000 : _GEN_268; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_270 = 9'h107 == addrEven[9:1] ? 32'h293f105 : _GEN_269; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_271 = 9'h108 == addrEven[9:1] ? 32'h400000 : _GEN_270; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_272 = 9'h109 == addrEven[9:1] ? 32'h3ff040 : _GEN_271; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_273 = 9'h10a == addrEven[9:1] ? 32'h87c20000 : _GEN_272; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_274 = 9'h10b == addrEven[9:1] ? 32'h87c40000 : _GEN_273; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_275 = 9'h10c == addrEven[9:1] ? 32'h2821100 : _GEN_274; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_276 = 9'h10d == addrEven[9:1] ? 32'h24c0030 : _GEN_275; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_277 = 9'h10e == addrEven[9:1] ? 32'hc800055 : _GEN_276; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_278 = 9'h10f == addrEven[9:1] ? 32'h20408 : _GEN_277; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_279 = 9'h110 == addrEven[9:1] ? 32'h400000 : _GEN_278; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_280 = 9'h111 == addrEven[9:1] ? 32'h2021466 : _GEN_279; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_281 = 9'h112 == addrEven[9:1] ? 32'h400000 : _GEN_280; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_282 = 9'h113 == addrEven[9:1] ? 32'h87c20000 : _GEN_281; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_283 = 9'h114 == addrEven[9:1] ? 32'h2821080 : _GEN_282; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_284 = 9'h115 == addrEven[9:1] ? 32'h1c21002 : _GEN_283; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_285 = 9'h116 == addrEven[9:1] ? 32'hcbffffa : _GEN_284; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_286 = 9'h117 == addrEven[9:1] ? 32'hf0080000 : _GEN_285; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_287 = 9'h118 == addrEven[9:1] ? 32'h87c40000 : _GEN_286; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_288 = 9'h119 == addrEven[9:1] ? 32'h87c21006 : _GEN_287; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_289 = 9'h11a == addrEven[9:1] ? 32'h2c42080 : _GEN_288; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_290 = 9'h11b == addrEven[9:1] ? 32'h87c20000 : _GEN_289; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_291 = 9'h11c == addrEven[9:1] ? 32'h2821080 : _GEN_290; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_292 = 9'h11d == addrEven[9:1] ? 32'h1c21002 : _GEN_291; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_293 = 9'h11e == addrEven[9:1] ? 32'hcbffffa : _GEN_292; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_294 = 9'h11f == addrEven[9:1] ? 32'h87c20000 : _GEN_293; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_295 = 9'h120 == addrEven[9:1] ? 32'hcc0000e : _GEN_294; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_296 = 9'h121 == addrEven[9:1] ? 32'h400000 : _GEN_295; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_297 = 9'h122 == addrEven[9:1] ? 32'h20000 : _GEN_296; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_298 = 9'h123 == addrEven[9:1] ? 32'h400000 : _GEN_297; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_299 = 9'h124 == addrEven[9:1] ? 32'h20004 : _GEN_298; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_300 = 9'h125 == addrEven[9:1] ? 32'h23001 : _GEN_299; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_301 = 9'h126 == addrEven[9:1] ? 32'h1c213ff : _GEN_300; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_302 = 9'h127 == addrEven[9:1] ? 32'h87c40000 : _GEN_301; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_303 = 9'h128 == addrEven[9:1] ? 32'h2842080 : _GEN_302; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_304 = 9'h129 == addrEven[9:1] ? 32'h1c42002 : _GEN_303; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_305 = 9'h12a == addrEven[9:1] ? 32'hcbffffa : _GEN_304; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_306 = 9'h12b == addrEven[9:1] ? 32'hf0080000 : _GEN_305; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_307 = 9'h12c == addrEven[9:1] ? 32'h400000 : _GEN_306; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_308 = 9'h12d == addrEven[9:1] ? 32'h1c42300 : _GEN_307; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_309 = 9'h12e == addrEven[9:1] ? 32'h87c40000 : _GEN_308; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_310 = 9'h12f == addrEven[9:1] ? 32'h2842100 : _GEN_309; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_311 = 9'h130 == addrEven[9:1] ? 32'h2063080 : _GEN_310; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_312 = 9'h131 == addrEven[9:1] ? 32'h1c813ff : _GEN_311; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_313 = 9'h132 == addrEven[9:1] ? 32'h20004 : _GEN_312; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_314 = 9'h133 == addrEven[9:1] ? 32'h87ca2000 : _GEN_313; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_315 = 9'h134 == addrEven[9:1] ? 32'h2d45200 : _GEN_314; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_316 = 9'h135 == addrEven[9:1] ? 32'h21001 : _GEN_315; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_317 = 9'h136 == addrEven[9:1] ? 32'h42001 : _GEN_316; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_318 = 9'h137 == addrEven[9:1] ? 32'h87c20000 : _GEN_317; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_319 = 9'h138 == addrEven[9:1] ? 32'h2c41100 : _GEN_318; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_320 = 9'h139 == addrEven[9:1] ? 32'h20404 : _GEN_319; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_321 = 9'h13a == addrEven[9:1] ? 32'h400000 : _GEN_320; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_322 = 9'h13b == addrEven[9:1] ? 32'h20004 : _GEN_321; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_323 = 9'h13c == addrEven[9:1] ? 32'h1c633ff : _GEN_322; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_324 = 9'h13d == addrEven[9:1] ? 32'h2821900 : _GEN_323; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_325 = 9'h13e == addrEven[9:1] ? 32'h2406020 : _GEN_324; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_326 = 9'h13f == addrEven[9:1] ? 32'h0 : _GEN_325; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_327 = 9'h140 == addrEven[9:1] ? 32'h0 : _GEN_326; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_328 = 9'h141 == addrEven[9:1] ? 32'h0 : _GEN_327; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_329 = 9'h142 == addrEven[9:1] ? 32'h0 : _GEN_328; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_330 = 9'h143 == addrEven[9:1] ? 32'h0 : _GEN_329; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_331 = 9'h144 == addrEven[9:1] ? 32'h0 : _GEN_330; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_332 = 9'h145 == addrEven[9:1] ? 32'h0 : _GEN_331; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_333 = 9'h146 == addrEven[9:1] ? 32'h0 : _GEN_332; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_334 = 9'h147 == addrEven[9:1] ? 32'h0 : _GEN_333; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_335 = 9'h148 == addrEven[9:1] ? 32'h0 : _GEN_334; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_336 = 9'h149 == addrEven[9:1] ? 32'h0 : _GEN_335; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_337 = 9'h14a == addrEven[9:1] ? 32'h0 : _GEN_336; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_338 = 9'h14b == addrEven[9:1] ? 32'h0 : _GEN_337; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_339 = 9'h14c == addrEven[9:1] ? 32'h0 : _GEN_338; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_340 = 9'h14d == addrEven[9:1] ? 32'h0 : _GEN_339; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_341 = 9'h14e == addrEven[9:1] ? 32'h0 : _GEN_340; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_342 = 9'h14f == addrEven[9:1] ? 32'h0 : _GEN_341; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_343 = 9'h150 == addrEven[9:1] ? 32'h0 : _GEN_342; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_344 = 9'h151 == addrEven[9:1] ? 32'h0 : _GEN_343; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_345 = 9'h152 == addrEven[9:1] ? 32'h0 : _GEN_344; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_346 = 9'h153 == addrEven[9:1] ? 32'h0 : _GEN_345; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_347 = 9'h154 == addrEven[9:1] ? 32'h0 : _GEN_346; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_348 = 9'h155 == addrEven[9:1] ? 32'h0 : _GEN_347; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_349 = 9'h156 == addrEven[9:1] ? 32'h0 : _GEN_348; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_350 = 9'h157 == addrEven[9:1] ? 32'h0 : _GEN_349; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_351 = 9'h158 == addrEven[9:1] ? 32'h0 : _GEN_350; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_352 = 9'h159 == addrEven[9:1] ? 32'h0 : _GEN_351; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_353 = 9'h15a == addrEven[9:1] ? 32'h0 : _GEN_352; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_354 = 9'h15b == addrEven[9:1] ? 32'h0 : _GEN_353; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_355 = 9'h15c == addrEven[9:1] ? 32'h0 : _GEN_354; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_356 = 9'h15d == addrEven[9:1] ? 32'h0 : _GEN_355; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_357 = 9'h15e == addrEven[9:1] ? 32'h0 : _GEN_356; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_358 = 9'h15f == addrEven[9:1] ? 32'h0 : _GEN_357; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_359 = 9'h160 == addrEven[9:1] ? 32'h0 : _GEN_358; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_360 = 9'h161 == addrEven[9:1] ? 32'h0 : _GEN_359; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_361 = 9'h162 == addrEven[9:1] ? 32'h0 : _GEN_360; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_362 = 9'h163 == addrEven[9:1] ? 32'h0 : _GEN_361; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_363 = 9'h164 == addrEven[9:1] ? 32'h0 : _GEN_362; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_364 = 9'h165 == addrEven[9:1] ? 32'h0 : _GEN_363; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_365 = 9'h166 == addrEven[9:1] ? 32'h0 : _GEN_364; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_366 = 9'h167 == addrEven[9:1] ? 32'h0 : _GEN_365; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_367 = 9'h168 == addrEven[9:1] ? 32'h0 : _GEN_366; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_368 = 9'h169 == addrEven[9:1] ? 32'h0 : _GEN_367; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_369 = 9'h16a == addrEven[9:1] ? 32'h0 : _GEN_368; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_370 = 9'h16b == addrEven[9:1] ? 32'h0 : _GEN_369; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_371 = 9'h16c == addrEven[9:1] ? 32'h0 : _GEN_370; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_372 = 9'h16d == addrEven[9:1] ? 32'h0 : _GEN_371; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_373 = 9'h16e == addrEven[9:1] ? 32'h0 : _GEN_372; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_374 = 9'h16f == addrEven[9:1] ? 32'h0 : _GEN_373; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_375 = 9'h170 == addrEven[9:1] ? 32'h0 : _GEN_374; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_376 = 9'h171 == addrEven[9:1] ? 32'h0 : _GEN_375; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_377 = 9'h172 == addrEven[9:1] ? 32'h0 : _GEN_376; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_378 = 9'h173 == addrEven[9:1] ? 32'h0 : _GEN_377; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_379 = 9'h174 == addrEven[9:1] ? 32'h0 : _GEN_378; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_380 = 9'h175 == addrEven[9:1] ? 32'h0 : _GEN_379; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_381 = 9'h176 == addrEven[9:1] ? 32'h0 : _GEN_380; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_382 = 9'h177 == addrEven[9:1] ? 32'h0 : _GEN_381; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_383 = 9'h178 == addrEven[9:1] ? 32'h0 : _GEN_382; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_384 = 9'h179 == addrEven[9:1] ? 32'h0 : _GEN_383; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_385 = 9'h17a == addrEven[9:1] ? 32'h0 : _GEN_384; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_386 = 9'h17b == addrEven[9:1] ? 32'h0 : _GEN_385; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_387 = 9'h17c == addrEven[9:1] ? 32'h0 : _GEN_386; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_388 = 9'h17d == addrEven[9:1] ? 32'h0 : _GEN_387; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_389 = 9'h17e == addrEven[9:1] ? 32'h0 : _GEN_388; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_390 = 9'h17f == addrEven[9:1] ? 32'h0 : _GEN_389; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_391 = 9'h180 == addrEven[9:1] ? 32'h0 : _GEN_390; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_392 = 9'h181 == addrEven[9:1] ? 32'h0 : _GEN_391; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_393 = 9'h182 == addrEven[9:1] ? 32'h0 : _GEN_392; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_394 = 9'h183 == addrEven[9:1] ? 32'h0 : _GEN_393; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_395 = 9'h184 == addrEven[9:1] ? 32'h0 : _GEN_394; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_396 = 9'h185 == addrEven[9:1] ? 32'h0 : _GEN_395; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_397 = 9'h186 == addrEven[9:1] ? 32'h0 : _GEN_396; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_398 = 9'h187 == addrEven[9:1] ? 32'h0 : _GEN_397; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_399 = 9'h188 == addrEven[9:1] ? 32'h0 : _GEN_398; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_400 = 9'h189 == addrEven[9:1] ? 32'h0 : _GEN_399; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_401 = 9'h18a == addrEven[9:1] ? 32'h0 : _GEN_400; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_402 = 9'h18b == addrEven[9:1] ? 32'h0 : _GEN_401; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_403 = 9'h18c == addrEven[9:1] ? 32'h0 : _GEN_402; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_404 = 9'h18d == addrEven[9:1] ? 32'h0 : _GEN_403; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_405 = 9'h18e == addrEven[9:1] ? 32'h0 : _GEN_404; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_406 = 9'h18f == addrEven[9:1] ? 32'h0 : _GEN_405; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_407 = 9'h190 == addrEven[9:1] ? 32'h0 : _GEN_406; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_408 = 9'h191 == addrEven[9:1] ? 32'h0 : _GEN_407; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_409 = 9'h192 == addrEven[9:1] ? 32'h0 : _GEN_408; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_410 = 9'h193 == addrEven[9:1] ? 32'h0 : _GEN_409; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_411 = 9'h194 == addrEven[9:1] ? 32'h0 : _GEN_410; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_412 = 9'h195 == addrEven[9:1] ? 32'h0 : _GEN_411; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_413 = 9'h196 == addrEven[9:1] ? 32'h0 : _GEN_412; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_414 = 9'h197 == addrEven[9:1] ? 32'h0 : _GEN_413; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_415 = 9'h198 == addrEven[9:1] ? 32'h0 : _GEN_414; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_416 = 9'h199 == addrEven[9:1] ? 32'h0 : _GEN_415; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_417 = 9'h19a == addrEven[9:1] ? 32'h0 : _GEN_416; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_418 = 9'h19b == addrEven[9:1] ? 32'h0 : _GEN_417; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_419 = 9'h19c == addrEven[9:1] ? 32'h0 : _GEN_418; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_420 = 9'h19d == addrEven[9:1] ? 32'h0 : _GEN_419; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_421 = 9'h19e == addrEven[9:1] ? 32'h0 : _GEN_420; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_422 = 9'h19f == addrEven[9:1] ? 32'h0 : _GEN_421; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_423 = 9'h1a0 == addrEven[9:1] ? 32'h0 : _GEN_422; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_424 = 9'h1a1 == addrEven[9:1] ? 32'h0 : _GEN_423; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_425 = 9'h1a2 == addrEven[9:1] ? 32'h0 : _GEN_424; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_426 = 9'h1a3 == addrEven[9:1] ? 32'h0 : _GEN_425; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_427 = 9'h1a4 == addrEven[9:1] ? 32'h0 : _GEN_426; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_428 = 9'h1a5 == addrEven[9:1] ? 32'h0 : _GEN_427; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_429 = 9'h1a6 == addrEven[9:1] ? 32'h0 : _GEN_428; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_430 = 9'h1a7 == addrEven[9:1] ? 32'h0 : _GEN_429; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_431 = 9'h1a8 == addrEven[9:1] ? 32'h0 : _GEN_430; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_432 = 9'h1a9 == addrEven[9:1] ? 32'h0 : _GEN_431; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_433 = 9'h1aa == addrEven[9:1] ? 32'h0 : _GEN_432; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_434 = 9'h1ab == addrEven[9:1] ? 32'h0 : _GEN_433; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_435 = 9'h1ac == addrEven[9:1] ? 32'h0 : _GEN_434; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_436 = 9'h1ad == addrEven[9:1] ? 32'h0 : _GEN_435; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_437 = 9'h1ae == addrEven[9:1] ? 32'h0 : _GEN_436; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_438 = 9'h1af == addrEven[9:1] ? 32'h0 : _GEN_437; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_439 = 9'h1b0 == addrEven[9:1] ? 32'h0 : _GEN_438; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_440 = 9'h1b1 == addrEven[9:1] ? 32'h0 : _GEN_439; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_441 = 9'h1b2 == addrEven[9:1] ? 32'h0 : _GEN_440; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_442 = 9'h1b3 == addrEven[9:1] ? 32'h0 : _GEN_441; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_443 = 9'h1b4 == addrEven[9:1] ? 32'h0 : _GEN_442; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_444 = 9'h1b5 == addrEven[9:1] ? 32'h0 : _GEN_443; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_445 = 9'h1b6 == addrEven[9:1] ? 32'h0 : _GEN_444; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_446 = 9'h1b7 == addrEven[9:1] ? 32'h0 : _GEN_445; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_447 = 9'h1b8 == addrEven[9:1] ? 32'h0 : _GEN_446; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_448 = 9'h1b9 == addrEven[9:1] ? 32'h0 : _GEN_447; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_449 = 9'h1ba == addrEven[9:1] ? 32'h0 : _GEN_448; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_450 = 9'h1bb == addrEven[9:1] ? 32'h0 : _GEN_449; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_451 = 9'h1bc == addrEven[9:1] ? 32'h0 : _GEN_450; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_452 = 9'h1bd == addrEven[9:1] ? 32'h0 : _GEN_451; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_453 = 9'h1be == addrEven[9:1] ? 32'h0 : _GEN_452; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_454 = 9'h1bf == addrEven[9:1] ? 32'h0 : _GEN_453; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_455 = 9'h1c0 == addrEven[9:1] ? 32'h0 : _GEN_454; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_456 = 9'h1c1 == addrEven[9:1] ? 32'h0 : _GEN_455; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_457 = 9'h1c2 == addrEven[9:1] ? 32'h0 : _GEN_456; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_458 = 9'h1c3 == addrEven[9:1] ? 32'h0 : _GEN_457; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_459 = 9'h1c4 == addrEven[9:1] ? 32'h0 : _GEN_458; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_460 = 9'h1c5 == addrEven[9:1] ? 32'h0 : _GEN_459; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_461 = 9'h1c6 == addrEven[9:1] ? 32'h0 : _GEN_460; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_462 = 9'h1c7 == addrEven[9:1] ? 32'h0 : _GEN_461; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_463 = 9'h1c8 == addrEven[9:1] ? 32'h0 : _GEN_462; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_464 = 9'h1c9 == addrEven[9:1] ? 32'h0 : _GEN_463; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_465 = 9'h1ca == addrEven[9:1] ? 32'h0 : _GEN_464; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_466 = 9'h1cb == addrEven[9:1] ? 32'h0 : _GEN_465; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_467 = 9'h1cc == addrEven[9:1] ? 32'h0 : _GEN_466; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_468 = 9'h1cd == addrEven[9:1] ? 32'h0 : _GEN_467; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_469 = 9'h1ce == addrEven[9:1] ? 32'h0 : _GEN_468; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_470 = 9'h1cf == addrEven[9:1] ? 32'h0 : _GEN_469; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_471 = 9'h1d0 == addrEven[9:1] ? 32'h0 : _GEN_470; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_472 = 9'h1d1 == addrEven[9:1] ? 32'h0 : _GEN_471; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_473 = 9'h1d2 == addrEven[9:1] ? 32'h0 : _GEN_472; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_474 = 9'h1d3 == addrEven[9:1] ? 32'h0 : _GEN_473; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_475 = 9'h1d4 == addrEven[9:1] ? 32'h0 : _GEN_474; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_476 = 9'h1d5 == addrEven[9:1] ? 32'h0 : _GEN_475; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_477 = 9'h1d6 == addrEven[9:1] ? 32'h0 : _GEN_476; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_478 = 9'h1d7 == addrEven[9:1] ? 32'h0 : _GEN_477; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_479 = 9'h1d8 == addrEven[9:1] ? 32'h0 : _GEN_478; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_480 = 9'h1d9 == addrEven[9:1] ? 32'h0 : _GEN_479; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_481 = 9'h1da == addrEven[9:1] ? 32'h0 : _GEN_480; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_482 = 9'h1db == addrEven[9:1] ? 32'h0 : _GEN_481; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_483 = 9'h1dc == addrEven[9:1] ? 32'h0 : _GEN_482; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_484 = 9'h1dd == addrEven[9:1] ? 32'h0 : _GEN_483; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_485 = 9'h1de == addrEven[9:1] ? 32'h0 : _GEN_484; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_486 = 9'h1df == addrEven[9:1] ? 32'h0 : _GEN_485; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_487 = 9'h1e0 == addrEven[9:1] ? 32'h0 : _GEN_486; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_488 = 9'h1e1 == addrEven[9:1] ? 32'h0 : _GEN_487; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_489 = 9'h1e2 == addrEven[9:1] ? 32'h0 : _GEN_488; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_490 = 9'h1e3 == addrEven[9:1] ? 32'h0 : _GEN_489; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_491 = 9'h1e4 == addrEven[9:1] ? 32'h0 : _GEN_490; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_492 = 9'h1e5 == addrEven[9:1] ? 32'h0 : _GEN_491; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_493 = 9'h1e6 == addrEven[9:1] ? 32'h0 : _GEN_492; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_494 = 9'h1e7 == addrEven[9:1] ? 32'h0 : _GEN_493; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_495 = 9'h1e8 == addrEven[9:1] ? 32'h0 : _GEN_494; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_496 = 9'h1e9 == addrEven[9:1] ? 32'h0 : _GEN_495; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_497 = 9'h1ea == addrEven[9:1] ? 32'h0 : _GEN_496; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_498 = 9'h1eb == addrEven[9:1] ? 32'h0 : _GEN_497; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_499 = 9'h1ec == addrEven[9:1] ? 32'h0 : _GEN_498; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_500 = 9'h1ed == addrEven[9:1] ? 32'h0 : _GEN_499; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_501 = 9'h1ee == addrEven[9:1] ? 32'h0 : _GEN_500; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_502 = 9'h1ef == addrEven[9:1] ? 32'h0 : _GEN_501; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_503 = 9'h1f0 == addrEven[9:1] ? 32'h0 : _GEN_502; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_504 = 9'h1f1 == addrEven[9:1] ? 32'h0 : _GEN_503; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_505 = 9'h1f2 == addrEven[9:1] ? 32'h0 : _GEN_504; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_506 = 9'h1f3 == addrEven[9:1] ? 32'h0 : _GEN_505; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_507 = 9'h1f4 == addrEven[9:1] ? 32'h0 : _GEN_506; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_508 = 9'h1f5 == addrEven[9:1] ? 32'h0 : _GEN_507; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_509 = 9'h1f6 == addrEven[9:1] ? 32'h0 : _GEN_508; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_510 = 9'h1f7 == addrEven[9:1] ? 32'h0 : _GEN_509; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_511 = 9'h1f8 == addrEven[9:1] ? 32'h0 : _GEN_510; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_512 = 9'h1f9 == addrEven[9:1] ? 32'h0 : _GEN_511; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_513 = 9'h1fa == addrEven[9:1] ? 32'h0 : _GEN_512; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_514 = 9'h1fb == addrEven[9:1] ? 32'h0 : _GEN_513; // @[Fetch.scala 100:26 Fetch.scala 100:26]
  wire [31:0] _GEN_520 = 9'h1 == addrOdd[9:1] ? 32'h87c40000 : 32'h87c20000; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_521 = 9'h2 == addrOdd[9:1] ? 32'h3e1000 : _GEN_520; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_522 = 9'h3 == addrOdd[9:1] ? 32'h2402026 : _GEN_521; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_523 = 9'h4 == addrOdd[9:1] ? 32'hf0010000 : _GEN_522; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_524 = 9'h5 == addrOdd[9:1] ? 32'h400000 : _GEN_523; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_525 = 9'h6 == addrOdd[9:1] ? 32'hcfc40000 : _GEN_524; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_526 = 9'h7 == addrOdd[9:1] ? 32'hcfc20000 : _GEN_525; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_527 = 9'h8 == addrOdd[9:1] ? 32'h4ac22085 : _GEN_526; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_528 = 9'h9 == addrOdd[9:1] ? 32'h400000 : _GEN_527; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_529 = 9'ha == addrOdd[9:1] ? 32'h4800000 : _GEN_528; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_530 = 9'hb == addrOdd[9:1] ? 32'h7ff024 : _GEN_529; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_531 = 9'hc == addrOdd[9:1] ? 32'h2c5f482 : _GEN_530; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_532 = 9'hd == addrOdd[9:1] ? 32'h2520037 : _GEN_531; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_533 = 9'he == addrOdd[9:1] ? 32'h2520030 : _GEN_532; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_534 = 9'hf == addrOdd[9:1] ? 32'h2c5fa83 : _GEN_533; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_535 = 9'h10 == addrOdd[9:1] ? 32'h2c5fb85 : _GEN_534; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_536 = 9'h11 == addrOdd[9:1] ? 32'h2c5fc87 : _GEN_535; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_537 = 9'h12 == addrOdd[9:1] ? 32'hf0020000 : _GEN_536; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_538 = 9'h13 == addrOdd[9:1] ? 32'h4403e8 : _GEN_537; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_539 = 9'h14 == addrOdd[9:1] ? 32'h87c40000 : _GEN_538; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_540 = 9'h15 == addrOdd[9:1] ? 32'h2842083 : _GEN_539; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_541 = 9'h16 == addrOdd[9:1] ? 32'h2041100 : _GEN_540; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_542 = 9'h17 == addrOdd[9:1] ? 32'hcbffffa : _GEN_541; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_543 = 9'h18 == addrOdd[9:1] ? 32'h2c60004 : _GEN_542; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_544 = 9'h19 == addrOdd[9:1] ? 32'hf0000000 : _GEN_543; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_545 = 9'h1a == addrOdd[9:1] ? 32'h400000 : _GEN_544; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_546 = 9'h1b == addrOdd[9:1] ? 32'h4c800023 : _GEN_545; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_547 = 9'h1c == addrOdd[9:1] ? 32'hf0000000 : _GEN_546; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_548 = 9'h1d == addrOdd[9:1] ? 32'h400000 : _GEN_547; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_549 = 9'h1e == addrOdd[9:1] ? 32'h2c62009 : _GEN_548; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_550 = 9'h1f == addrOdd[9:1] ? 32'h460001 : _GEN_549; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_551 = 9'h20 == addrOdd[9:1] ? 32'h2c62188 : _GEN_550; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_552 = 9'h21 == addrOdd[9:1] ? 32'h400000 : _GEN_551; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_553 = 9'h22 == addrOdd[9:1] ? 32'h2c62007 : _GEN_552; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_554 = 9'h23 == addrOdd[9:1] ? 32'h400000 : _GEN_553; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_555 = 9'h24 == addrOdd[9:1] ? 32'h2c61006 : _GEN_554; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_556 = 9'h25 == addrOdd[9:1] ? 32'h87c20000 : _GEN_555; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_557 = 9'h26 == addrOdd[9:1] ? 32'h2821080 : _GEN_556; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_558 = 9'h27 == addrOdd[9:1] ? 32'hc21004 : _GEN_557; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_559 = 9'h28 == addrOdd[9:1] ? 32'h2820185 : _GEN_558; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_560 = 9'h29 == addrOdd[9:1] ? 32'h20210e1 : _GEN_559; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_561 = 9'h2a == addrOdd[9:1] ? 32'h2820185 : _GEN_560; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_562 = 9'h2b == addrOdd[9:1] ? 32'h2021161 : _GEN_561; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_563 = 9'h2c == addrOdd[9:1] ? 32'h480001d : _GEN_562; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_564 = 9'h2d == addrOdd[9:1] ? 32'hf0000000 : _GEN_563; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_565 = 9'h2e == addrOdd[9:1] ? 32'h400000 : _GEN_564; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_566 = 9'h2f == addrOdd[9:1] ? 32'hcc00010 : _GEN_565; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_567 = 9'h30 == addrOdd[9:1] ? 32'h40000 : _GEN_566; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_568 = 9'h31 == addrOdd[9:1] ? 32'h2c61009 : _GEN_567; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_569 = 9'h32 == addrOdd[9:1] ? 32'h2c61188 : _GEN_568; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_570 = 9'h33 == addrOdd[9:1] ? 32'h2c61006 : _GEN_569; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_571 = 9'h34 == addrOdd[9:1] ? 32'h87c60000 : _GEN_570; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_572 = 9'h35 == addrOdd[9:1] ? 32'h2863082 : _GEN_571; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_573 = 9'h36 == addrOdd[9:1] ? 32'h20221b4 : _GEN_572; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_574 = 9'h37 == addrOdd[9:1] ? 32'h421001 : _GEN_573; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_575 = 9'h38 == addrOdd[9:1] ? 32'hcfffffe : _GEN_574; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_576 = 9'h39 == addrOdd[9:1] ? 32'h2c60105 : _GEN_575; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_577 = 9'h3a == addrOdd[9:1] ? 32'h2c60084 : _GEN_576; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_578 = 9'h3b == addrOdd[9:1] ? 32'hf0000000 : _GEN_577; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_579 = 9'h3c == addrOdd[9:1] ? 32'h400000 : _GEN_578; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_580 = 9'h3d == addrOdd[9:1] ? 32'h20000 : _GEN_579; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_581 = 9'h3e == addrOdd[9:1] ? 32'h87c4100d : _GEN_580; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_582 = 9'h3f == addrOdd[9:1] ? 32'h2862180 : _GEN_581; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_583 = 9'h40 == addrOdd[9:1] ? 32'h2c22180 : _GEN_582; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_584 = 9'h41 == addrOdd[9:1] ? 32'hf0000000 : _GEN_583; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_585 = 9'h42 == addrOdd[9:1] ? 32'h21001 : _GEN_584; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_586 = 9'h43 == addrOdd[9:1] ? 32'h2021134 : _GEN_585; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_587 = 9'h44 == addrOdd[9:1] ? 32'h87c20000 : _GEN_586; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_588 = 9'h45 == addrOdd[9:1] ? 32'h2821080 : _GEN_587; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_589 = 9'h46 == addrOdd[9:1] ? 32'h2021031 : _GEN_588; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_590 = 9'h47 == addrOdd[9:1] ? 32'h87c20000 : _GEN_589; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_591 = 9'h48 == addrOdd[9:1] ? 32'h2821080 : _GEN_590; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_592 = 9'h49 == addrOdd[9:1] ? 32'h4c00016 : _GEN_591; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_593 = 9'h4a == addrOdd[9:1] ? 32'h2c61109 : _GEN_592; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_594 = 9'h4b == addrOdd[9:1] ? 32'h2c60085 : _GEN_593; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_595 = 9'h4c == addrOdd[9:1] ? 32'hf0000000 : _GEN_594; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_596 = 9'h4d == addrOdd[9:1] ? 32'h20001 : _GEN_595; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_597 = 9'h4e == addrOdd[9:1] ? 32'hc80000c : _GEN_596; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_598 = 9'h4f == addrOdd[9:1] ? 32'h2842189 : _GEN_597; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_599 = 9'h50 == addrOdd[9:1] ? 32'h2022161 : _GEN_598; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_600 = 9'h51 == addrOdd[9:1] ? 32'h87c40000 : _GEN_599; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_601 = 9'h52 == addrOdd[9:1] ? 32'h2842082 : _GEN_600; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_602 = 9'h53 == addrOdd[9:1] ? 32'h2021134 : _GEN_601; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_603 = 9'h54 == addrOdd[9:1] ? 32'h2840184 : _GEN_602; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_604 = 9'h55 == addrOdd[9:1] ? 32'h2022060 : _GEN_603; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_605 = 9'h56 == addrOdd[9:1] ? 32'h87c20000 : _GEN_604; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_606 = 9'h57 == addrOdd[9:1] ? 32'h2821085 : _GEN_605; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_607 = 9'h58 == addrOdd[9:1] ? 32'h20220b2 : _GEN_606; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_608 = 9'h59 == addrOdd[9:1] ? 32'hf0010000 : _GEN_607; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_609 = 9'h5a == addrOdd[9:1] ? 32'h80000000 : _GEN_608; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_610 = 9'h5b == addrOdd[9:1] ? 32'h400000 : _GEN_609; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_611 = 9'h5c == addrOdd[9:1] ? 32'h2820184 : _GEN_610; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_612 = 9'h5d == addrOdd[9:1] ? 32'h6001004 : _GEN_611; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_613 = 9'h5e == addrOdd[9:1] ? 32'hf0010000 : _GEN_612; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_614 = 9'h5f == addrOdd[9:1] ? 32'h400000 : _GEN_613; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_615 = 9'h60 == addrOdd[9:1] ? 32'hcfc60000 : _GEN_614; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_616 = 9'h61 == addrOdd[9:1] ? 32'hcfc40000 : _GEN_615; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_617 = 9'h62 == addrOdd[9:1] ? 32'h4ac23105 : _GEN_616; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_618 = 9'h63 == addrOdd[9:1] ? 32'h400000 : _GEN_617; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_619 = 9'h64 == addrOdd[9:1] ? 32'hf0000000 : _GEN_618; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_620 = 9'h65 == addrOdd[9:1] ? 32'h400000 : _GEN_619; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_621 = 9'h66 == addrOdd[9:1] ? 32'h2c62088 : _GEN_620; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_622 = 9'h67 == addrOdd[9:1] ? 32'h87c40000 : _GEN_621; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_623 = 9'h68 == addrOdd[9:1] ? 32'h2842080 : _GEN_622; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_624 = 9'h69 == addrOdd[9:1] ? 32'h2022031 : _GEN_623; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_625 = 9'h6a == addrOdd[9:1] ? 32'h40004 : _GEN_624; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_626 = 9'h6b == addrOdd[9:1] ? 32'hf0000000 : _GEN_625; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_627 = 9'h6c == addrOdd[9:1] ? 32'h400000 : _GEN_626; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_628 = 9'h6d == addrOdd[9:1] ? 32'h2c61109 : _GEN_627; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_629 = 9'h6e == addrOdd[9:1] ? 32'h400000 : _GEN_628; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_630 = 9'h6f == addrOdd[9:1] ? 32'hcbffff7 : _GEN_629; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_631 = 9'h70 == addrOdd[9:1] ? 32'hf0000000 : _GEN_630; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_632 = 9'h71 == addrOdd[9:1] ? 32'h4c00048 : _GEN_631; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_633 = 9'h72 == addrOdd[9:1] ? 32'h2c61009 : _GEN_632; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_634 = 9'h73 == addrOdd[9:1] ? 32'hf0000000 : _GEN_633; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_635 = 9'h74 == addrOdd[9:1] ? 32'h40001 : _GEN_634; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_636 = 9'h75 == addrOdd[9:1] ? 32'hc800011 : _GEN_635; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_637 = 9'h76 == addrOdd[9:1] ? 32'h2863189 : _GEN_636; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_638 = 9'h77 == addrOdd[9:1] ? 32'h2023060 : _GEN_637; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_639 = 9'h78 == addrOdd[9:1] ? 32'hc62004 : _GEN_638; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_640 = 9'h79 == addrOdd[9:1] ? 32'h400000 : _GEN_639; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_641 = 9'h7a == addrOdd[9:1] ? 32'hcbffffc : _GEN_640; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_642 = 9'h7b == addrOdd[9:1] ? 32'hf0000000 : _GEN_641; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_643 = 9'h7c == addrOdd[9:1] ? 32'h42001 : _GEN_642; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_644 = 9'h7d == addrOdd[9:1] ? 32'hcbffff1 : _GEN_643; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_645 = 9'h7e == addrOdd[9:1] ? 32'hf0080000 : _GEN_644; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_646 = 9'h7f == addrOdd[9:1] ? 32'h400000 : _GEN_645; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_647 = 9'h80 == addrOdd[9:1] ? 32'h4cbffffb : _GEN_646; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_648 = 9'h81 == addrOdd[9:1] ? 32'hf0080000 : _GEN_647; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_649 = 9'h82 == addrOdd[9:1] ? 32'h87c40000 : _GEN_648; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_650 = 9'h83 == addrOdd[9:1] ? 32'h2842080 : _GEN_649; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_651 = 9'h84 == addrOdd[9:1] ? 32'h2022036 : _GEN_650; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_652 = 9'h85 == addrOdd[9:1] ? 32'h40078 : _GEN_651; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_653 = 9'h86 == addrOdd[9:1] ? 32'hf0080000 : _GEN_652; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_654 = 9'h87 == addrOdd[9:1] ? 32'h87c40000 : _GEN_653; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_655 = 9'h88 == addrOdd[9:1] ? 32'h2842080 : _GEN_654; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_656 = 9'h89 == addrOdd[9:1] ? 32'h2022036 : _GEN_655; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_657 = 9'h8a == addrOdd[9:1] ? 32'h87c40000 : _GEN_656; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_658 = 9'h8b == addrOdd[9:1] ? 32'h2c22081 : _GEN_657; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_659 = 9'h8c == addrOdd[9:1] ? 32'h2c60085 : _GEN_658; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_660 = 9'h8d == addrOdd[9:1] ? 32'hf0000000 : _GEN_659; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_661 = 9'h8e == addrOdd[9:1] ? 32'h20001 : _GEN_660; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_662 = 9'h8f == addrOdd[9:1] ? 32'hc80000c : _GEN_661; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_663 = 9'h90 == addrOdd[9:1] ? 32'h2842189 : _GEN_662; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_664 = 9'h91 == addrOdd[9:1] ? 32'h2022260 : _GEN_663; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_665 = 9'h92 == addrOdd[9:1] ? 32'h87c40000 : _GEN_664; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_666 = 9'h93 == addrOdd[9:1] ? 32'h2842082 : _GEN_665; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_667 = 9'h94 == addrOdd[9:1] ? 32'h2021134 : _GEN_666; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_668 = 9'h95 == addrOdd[9:1] ? 32'h87c40000 : _GEN_667; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_669 = 9'h96 == addrOdd[9:1] ? 32'h20001 : _GEN_668; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_670 = 9'h97 == addrOdd[9:1] ? 32'h2c22085 : _GEN_669; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_671 = 9'h98 == addrOdd[9:1] ? 32'h2c22085 : _GEN_670; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_672 = 9'h99 == addrOdd[9:1] ? 32'h2aff105 : _GEN_671; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_673 = 9'h9a == addrOdd[9:1] ? 32'h2b3f107 : _GEN_672; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_674 = 9'h9b == addrOdd[9:1] ? 32'h293f102 : _GEN_673; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_675 = 9'h9c == addrOdd[9:1] ? 32'h2409028 : _GEN_674; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_676 = 9'h9d == addrOdd[9:1] ? 32'h400000 : _GEN_675; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_677 = 9'h9e == addrOdd[9:1] ? 32'h293f100 : _GEN_676; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_678 = 9'h9f == addrOdd[9:1] ? 32'h20000 : _GEN_677; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_679 = 9'ha0 == addrOdd[9:1] ? 32'h3ff024 : _GEN_678; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_680 = 9'ha1 == addrOdd[9:1] ? 32'h7ff040 : _GEN_679; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_681 = 9'ha2 == addrOdd[9:1] ? 32'h2c5f487 : _GEN_680; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_682 = 9'ha3 == addrOdd[9:1] ? 32'h20000 : _GEN_681; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_683 = 9'ha4 == addrOdd[9:1] ? 32'h2c5fe0f : _GEN_682; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_684 = 9'ha5 == addrOdd[9:1] ? 32'h2c5f486 : _GEN_683; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_685 = 9'ha6 == addrOdd[9:1] ? 32'h2c5f485 : _GEN_684; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_686 = 9'ha7 == addrOdd[9:1] ? 32'h2c5fb09 : _GEN_685; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_687 = 9'ha8 == addrOdd[9:1] ? 32'h2c5fc0b : _GEN_686; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_688 = 9'ha9 == addrOdd[9:1] ? 32'h2c5fd0d : _GEN_687; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_689 = 9'haa == addrOdd[9:1] ? 32'h20000 : _GEN_688; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_690 = 9'hab == addrOdd[9:1] ? 32'h20004 : _GEN_689; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_691 = 9'hac == addrOdd[9:1] ? 32'h2d41100 : _GEN_690; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_692 = 9'had == addrOdd[9:1] ? 32'h20000 : _GEN_691; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_693 = 9'hae == addrOdd[9:1] ? 32'h400000 : _GEN_692; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_694 = 9'haf == addrOdd[9:1] ? 32'h2c42080 : _GEN_693; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_695 = 9'hb0 == addrOdd[9:1] ? 32'h2021134 : _GEN_694; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_696 = 9'hb1 == addrOdd[9:1] ? 32'h87c40000 : _GEN_695; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_697 = 9'hb2 == addrOdd[9:1] ? 32'h2c42080 : _GEN_696; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_698 = 9'hb3 == addrOdd[9:1] ? 32'h80000 : _GEN_697; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_699 = 9'hb4 == addrOdd[9:1] ? 32'h2c5f003 : _GEN_698; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_700 = 9'hb5 == addrOdd[9:1] ? 32'h340000 : _GEN_699; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_701 = 9'hb6 == addrOdd[9:1] ? 32'h2c5f002 : _GEN_700; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_702 = 9'hb7 == addrOdd[9:1] ? 32'h2c5f001 : _GEN_701; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_703 = 9'hb8 == addrOdd[9:1] ? 32'h20408 : _GEN_702; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_704 = 9'hb9 == addrOdd[9:1] ? 32'h420001 : _GEN_703; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_705 = 9'hba == addrOdd[9:1] ? 32'h40000 : _GEN_704; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_706 = 9'hbb == addrOdd[9:1] ? 32'h381000 : _GEN_705; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_707 = 9'hbc == addrOdd[9:1] ? 32'h2e3000 : _GEN_706; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_708 = 9'hbd == addrOdd[9:1] ? 32'h87c20000 : _GEN_707; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_709 = 9'hbe == addrOdd[9:1] ? 32'h2c21d80 : _GEN_708; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_710 = 9'hbf == addrOdd[9:1] ? 32'h440001 : _GEN_709; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_711 = 9'hc0 == addrOdd[9:1] ? 32'hcfffff6 : _GEN_710; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_712 = 9'hc1 == addrOdd[9:1] ? 32'h60000 : _GEN_711; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_713 = 9'hc2 == addrOdd[9:1] ? 32'h2022b34 : _GEN_712; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_714 = 9'hc3 == addrOdd[9:1] ? 32'hc57008 : _GEN_713; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_715 = 9'hc4 == addrOdd[9:1] ? 32'h2061106 : _GEN_714; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_716 = 9'hc5 == addrOdd[9:1] ? 32'h5c004 : _GEN_715; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_717 = 9'hc6 == addrOdd[9:1] ? 32'hc800025 : _GEN_716; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_718 = 9'hc7 == addrOdd[9:1] ? 32'h60008 : _GEN_717; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_719 = 9'hc8 == addrOdd[9:1] ? 32'h2024036 : _GEN_718; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_720 = 9'hc9 == addrOdd[9:1] ? 32'hedb88320 : _GEN_719; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_721 = 9'hca == addrOdd[9:1] ? 32'h9044001 : _GEN_720; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_722 = 9'hcb == addrOdd[9:1] ? 32'h463001 : _GEN_721; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_723 = 9'hcc == addrOdd[9:1] ? 32'hcbffff7 : _GEN_722; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_724 = 9'hcd == addrOdd[9:1] ? 32'h206300b : _GEN_723; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_725 = 9'hce == addrOdd[9:1] ? 32'h28bf103 : _GEN_724; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_726 = 9'hcf == addrOdd[9:1] ? 32'h20a1286 : _GEN_725; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_727 = 9'hd0 == addrOdd[9:1] ? 32'h2021db4 : _GEN_726; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_728 = 9'hd1 == addrOdd[9:1] ? 32'h289f102 : _GEN_727; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_729 = 9'hd2 == addrOdd[9:1] ? 32'h2023261 : _GEN_728; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_730 = 9'hd3 == addrOdd[9:1] ? 32'h20004 : _GEN_729; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_731 = 9'hd4 == addrOdd[9:1] ? 32'hc800018 : _GEN_730; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_732 = 9'hd5 == addrOdd[9:1] ? 32'hf0008010 : _GEN_731; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_733 = 9'hd6 == addrOdd[9:1] ? 32'h25000 : _GEN_732; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_734 = 9'hd7 == addrOdd[9:1] ? 32'h4c00012 : _GEN_733; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_735 = 9'hd8 == addrOdd[9:1] ? 32'h2c5f284 : _GEN_734; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_736 = 9'hd9 == addrOdd[9:1] ? 32'h59000 : _GEN_735; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_737 = 9'hda == addrOdd[9:1] ? 32'h2035c00 : _GEN_736; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_738 = 9'hdb == addrOdd[9:1] ? 32'hfffffffc : _GEN_737; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_739 = 9'hdc == addrOdd[9:1] ? 32'h4c0000c : _GEN_738; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_740 = 9'hdd == addrOdd[9:1] ? 32'h400000 : _GEN_739; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_741 = 9'hde == addrOdd[9:1] ? 32'h4800004 : _GEN_740; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_742 = 9'hdf == addrOdd[9:1] ? 32'h4800002 : _GEN_741; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_743 = 9'he0 == addrOdd[9:1] ? 32'h283f101 : _GEN_742; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_744 = 9'he1 == addrOdd[9:1] ? 32'h37b001 : _GEN_743; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_745 = 9'he2 == addrOdd[9:1] ? 32'h2023230 : _GEN_744; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_746 = 9'he3 == addrOdd[9:1] ? 32'h20220c7 : _GEN_745; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_747 = 9'he4 == addrOdd[9:1] ? 32'h64003 : _GEN_746; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_748 = 9'he5 == addrOdd[9:1] ? 32'hfffffffc : _GEN_747; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_749 = 9'he6 == addrOdd[9:1] ? 32'hcc0000a : _GEN_748; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_750 = 9'he7 == addrOdd[9:1] ? 32'h2c5f202 : _GEN_749; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_751 = 9'he8 == addrOdd[9:1] ? 32'h63004 : _GEN_750; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_752 = 9'he9 == addrOdd[9:1] ? 32'hcfffffd : _GEN_751; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_753 = 9'hea == addrOdd[9:1] ? 32'hfffffffc : _GEN_752; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_754 = 9'heb == addrOdd[9:1] ? 32'h360002 : _GEN_753; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_755 = 9'hec == addrOdd[9:1] ? 32'h287f100 : _GEN_754; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_756 = 9'hed == addrOdd[9:1] ? 32'h63001 : _GEN_755; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_757 = 9'hee == addrOdd[9:1] ? 32'h2c5f202 : _GEN_756; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_758 = 9'hef == addrOdd[9:1] ? 32'h1c75003 : _GEN_757; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_759 = 9'hf0 == addrOdd[9:1] ? 32'h80a0000 : _GEN_758; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_760 = 9'hf1 == addrOdd[9:1] ? 32'h2c5f081 : _GEN_759; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_761 = 9'hf2 == addrOdd[9:1] ? 32'h3c003 : _GEN_760; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_762 = 9'hf3 == addrOdd[9:1] ? 32'hcffff90 : _GEN_761; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_763 = 9'hf4 == addrOdd[9:1] ? 32'h3c000 : _GEN_762; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_764 = 9'hf5 == addrOdd[9:1] ? 32'hf0080000 : _GEN_763; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_765 = 9'hf6 == addrOdd[9:1] ? 32'h400000 : _GEN_764; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_766 = 9'hf7 == addrOdd[9:1] ? 32'h4cbffffb : _GEN_765; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_767 = 9'hf8 == addrOdd[9:1] ? 32'h1c410ff : _GEN_766; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_768 = 9'hf9 == addrOdd[9:1] ? 32'hf0080000 : _GEN_767; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_769 = 9'hfa == addrOdd[9:1] ? 32'hcc0000c : _GEN_768; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_770 = 9'hfb == addrOdd[9:1] ? 32'h20000 : _GEN_769; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_771 = 9'hfc == addrOdd[9:1] ? 32'h285f104 : _GEN_770; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_772 = 9'hfd == addrOdd[9:1] ? 32'h2021131 : _GEN_771; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_773 = 9'hfe == addrOdd[9:1] ? 32'h20000 : _GEN_772; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_774 = 9'hff == addrOdd[9:1] ? 32'h283f101 : _GEN_773; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_775 = 9'h100 == addrOdd[9:1] ? 32'h2adf109 : _GEN_774; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_776 = 9'h101 == addrOdd[9:1] ? 32'h2b1f10b : _GEN_775; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_777 = 9'h102 == addrOdd[9:1] ? 32'h2b5f10d : _GEN_776; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_778 = 9'h103 == addrOdd[9:1] ? 32'h2b9f10f : _GEN_777; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_779 = 9'h104 == addrOdd[9:1] ? 32'h2abf108 : _GEN_778; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_780 = 9'h105 == addrOdd[9:1] ? 32'h293f106 : _GEN_779; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_781 = 9'h106 == addrOdd[9:1] ? 32'h2409027 : _GEN_780; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_782 = 9'h107 == addrOdd[9:1] ? 32'h6400000 : _GEN_781; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_783 = 9'h108 == addrOdd[9:1] ? 32'h2409020 : _GEN_782; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_784 = 9'h109 == addrOdd[9:1] ? 32'h1a4 : _GEN_783; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_785 = 9'h10a == addrOdd[9:1] ? 32'h20000 : _GEN_784; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_786 = 9'h10b == addrOdd[9:1] ? 32'h20404 : _GEN_785; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_787 = 9'h10c == addrOdd[9:1] ? 32'h2842100 : _GEN_786; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_788 = 9'h10d == addrOdd[9:1] ? 32'h20220b1 : _GEN_787; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_789 = 9'h10e == addrOdd[9:1] ? 32'h87c40000 : _GEN_788; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_790 = 9'h10f == addrOdd[9:1] ? 32'h2822100 : _GEN_789; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_791 = 9'h110 == addrOdd[9:1] ? 32'h1021001 : _GEN_790; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_792 = 9'h111 == addrOdd[9:1] ? 32'hcc00012 : _GEN_791; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_793 = 9'h112 == addrOdd[9:1] ? 32'h2c42080 : _GEN_792; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_794 = 9'h113 == addrOdd[9:1] ? 32'hf0080000 : _GEN_793; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_795 = 9'h114 == addrOdd[9:1] ? 32'h400000 : _GEN_794; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_796 = 9'h115 == addrOdd[9:1] ? 32'h2021060 : _GEN_795; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_797 = 9'h116 == addrOdd[9:1] ? 32'h87c20000 : _GEN_796; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_798 = 9'h117 == addrOdd[9:1] ? 32'h2821081 : _GEN_797; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_799 = 9'h118 == addrOdd[9:1] ? 32'h20408 : _GEN_798; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_800 = 9'h119 == addrOdd[9:1] ? 32'hff00 : _GEN_799; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_801 = 9'h11a == addrOdd[9:1] ? 32'h1c41001 : _GEN_800; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_802 = 9'h11b == addrOdd[9:1] ? 32'hf0080000 : _GEN_801; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_803 = 9'h11c == addrOdd[9:1] ? 32'h400000 : _GEN_802; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_804 = 9'h11d == addrOdd[9:1] ? 32'h2021060 : _GEN_803; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_805 = 9'h11e == addrOdd[9:1] ? 32'h2022060 : _GEN_804; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_806 = 9'h11f == addrOdd[9:1] ? 32'hf0080000 : _GEN_805; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_807 = 9'h120 == addrOdd[9:1] ? 32'h2821081 : _GEN_806; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_808 = 9'h121 == addrOdd[9:1] ? 32'h87c40000 : _GEN_807; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_809 = 9'h122 == addrOdd[9:1] ? 32'h2862100 : _GEN_808; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_810 = 9'h123 == addrOdd[9:1] ? 32'h87c83000 : _GEN_809; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_811 = 9'h124 == addrOdd[9:1] ? 32'h2d44080 : _GEN_810; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_812 = 9'h125 == addrOdd[9:1] ? 32'h4c00026 : _GEN_811; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_813 = 9'h126 == addrOdd[9:1] ? 32'h2c42080 : _GEN_812; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_814 = 9'h127 == addrOdd[9:1] ? 32'hf0080000 : _GEN_813; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_815 = 9'h128 == addrOdd[9:1] ? 32'h400000 : _GEN_814; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_816 = 9'h129 == addrOdd[9:1] ? 32'h2022060 : _GEN_815; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_817 = 9'h12a == addrOdd[9:1] ? 32'h87c40000 : _GEN_816; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_818 = 9'h12b == addrOdd[9:1] ? 32'h2862081 : _GEN_817; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_819 = 9'h12c == addrOdd[9:1] ? 32'hc43002 : _GEN_818; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_820 = 9'h12d == addrOdd[9:1] ? 32'h2022086 : _GEN_819; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_821 = 9'h12e == addrOdd[9:1] ? 32'h20000 : _GEN_820; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_822 = 9'h12f == addrOdd[9:1] ? 32'h1c6303f : _GEN_821; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_823 = 9'h130 == addrOdd[9:1] ? 32'h63002 : _GEN_822; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_824 = 9'h131 == addrOdd[9:1] ? 32'h87c84000 : _GEN_823; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_825 = 9'h132 == addrOdd[9:1] ? 32'h2884900 : _GEN_824; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_826 = 9'h133 == addrOdd[9:1] ? 32'h20004 : _GEN_825; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_827 = 9'h134 == addrOdd[9:1] ? 32'h20211b2 : _GEN_826; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_828 = 9'h135 == addrOdd[9:1] ? 32'hcfffff7 : _GEN_827; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_829 = 9'h136 == addrOdd[9:1] ? 32'h1c423ff : _GEN_828; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_830 = 9'h137 == addrOdd[9:1] ? 32'h20000 : _GEN_829; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_831 = 9'h138 == addrOdd[9:1] ? 32'h87c40000 : _GEN_830; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_832 = 9'h139 == addrOdd[9:1] ? 32'h2862100 : _GEN_831; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_833 = 9'h13a == addrOdd[9:1] ? 32'h87c23000 : _GEN_832; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_834 = 9'h13b == addrOdd[9:1] ? 32'h63001 : _GEN_833; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_835 = 9'h13c == addrOdd[9:1] ? 32'h6400000 : _GEN_834; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_836 = 9'h13d == addrOdd[9:1] ? 32'h2c42180 : _GEN_835; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_837 = 9'h13e == addrOdd[9:1] ? 32'h0 : _GEN_836; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_838 = 9'h13f == addrOdd[9:1] ? 32'h0 : _GEN_837; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_839 = 9'h140 == addrOdd[9:1] ? 32'h0 : _GEN_838; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_840 = 9'h141 == addrOdd[9:1] ? 32'h0 : _GEN_839; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_841 = 9'h142 == addrOdd[9:1] ? 32'h0 : _GEN_840; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_842 = 9'h143 == addrOdd[9:1] ? 32'h0 : _GEN_841; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_843 = 9'h144 == addrOdd[9:1] ? 32'h0 : _GEN_842; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_844 = 9'h145 == addrOdd[9:1] ? 32'h0 : _GEN_843; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_845 = 9'h146 == addrOdd[9:1] ? 32'h0 : _GEN_844; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_846 = 9'h147 == addrOdd[9:1] ? 32'h0 : _GEN_845; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_847 = 9'h148 == addrOdd[9:1] ? 32'h0 : _GEN_846; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_848 = 9'h149 == addrOdd[9:1] ? 32'h0 : _GEN_847; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_849 = 9'h14a == addrOdd[9:1] ? 32'h0 : _GEN_848; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_850 = 9'h14b == addrOdd[9:1] ? 32'h0 : _GEN_849; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_851 = 9'h14c == addrOdd[9:1] ? 32'h0 : _GEN_850; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_852 = 9'h14d == addrOdd[9:1] ? 32'h0 : _GEN_851; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_853 = 9'h14e == addrOdd[9:1] ? 32'h0 : _GEN_852; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_854 = 9'h14f == addrOdd[9:1] ? 32'h0 : _GEN_853; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_855 = 9'h150 == addrOdd[9:1] ? 32'h0 : _GEN_854; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_856 = 9'h151 == addrOdd[9:1] ? 32'h0 : _GEN_855; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_857 = 9'h152 == addrOdd[9:1] ? 32'h0 : _GEN_856; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_858 = 9'h153 == addrOdd[9:1] ? 32'h0 : _GEN_857; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_859 = 9'h154 == addrOdd[9:1] ? 32'h0 : _GEN_858; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_860 = 9'h155 == addrOdd[9:1] ? 32'h0 : _GEN_859; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_861 = 9'h156 == addrOdd[9:1] ? 32'h0 : _GEN_860; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_862 = 9'h157 == addrOdd[9:1] ? 32'h0 : _GEN_861; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_863 = 9'h158 == addrOdd[9:1] ? 32'h0 : _GEN_862; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_864 = 9'h159 == addrOdd[9:1] ? 32'h0 : _GEN_863; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_865 = 9'h15a == addrOdd[9:1] ? 32'h0 : _GEN_864; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_866 = 9'h15b == addrOdd[9:1] ? 32'h0 : _GEN_865; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_867 = 9'h15c == addrOdd[9:1] ? 32'h0 : _GEN_866; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_868 = 9'h15d == addrOdd[9:1] ? 32'h0 : _GEN_867; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_869 = 9'h15e == addrOdd[9:1] ? 32'h0 : _GEN_868; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_870 = 9'h15f == addrOdd[9:1] ? 32'h0 : _GEN_869; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_871 = 9'h160 == addrOdd[9:1] ? 32'h0 : _GEN_870; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_872 = 9'h161 == addrOdd[9:1] ? 32'h0 : _GEN_871; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_873 = 9'h162 == addrOdd[9:1] ? 32'h0 : _GEN_872; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_874 = 9'h163 == addrOdd[9:1] ? 32'h0 : _GEN_873; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_875 = 9'h164 == addrOdd[9:1] ? 32'h0 : _GEN_874; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_876 = 9'h165 == addrOdd[9:1] ? 32'h0 : _GEN_875; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_877 = 9'h166 == addrOdd[9:1] ? 32'h0 : _GEN_876; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_878 = 9'h167 == addrOdd[9:1] ? 32'h0 : _GEN_877; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_879 = 9'h168 == addrOdd[9:1] ? 32'h0 : _GEN_878; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_880 = 9'h169 == addrOdd[9:1] ? 32'h0 : _GEN_879; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_881 = 9'h16a == addrOdd[9:1] ? 32'h0 : _GEN_880; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_882 = 9'h16b == addrOdd[9:1] ? 32'h0 : _GEN_881; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_883 = 9'h16c == addrOdd[9:1] ? 32'h0 : _GEN_882; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_884 = 9'h16d == addrOdd[9:1] ? 32'h0 : _GEN_883; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_885 = 9'h16e == addrOdd[9:1] ? 32'h0 : _GEN_884; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_886 = 9'h16f == addrOdd[9:1] ? 32'h0 : _GEN_885; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_887 = 9'h170 == addrOdd[9:1] ? 32'h0 : _GEN_886; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_888 = 9'h171 == addrOdd[9:1] ? 32'h0 : _GEN_887; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_889 = 9'h172 == addrOdd[9:1] ? 32'h0 : _GEN_888; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_890 = 9'h173 == addrOdd[9:1] ? 32'h0 : _GEN_889; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_891 = 9'h174 == addrOdd[9:1] ? 32'h0 : _GEN_890; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_892 = 9'h175 == addrOdd[9:1] ? 32'h0 : _GEN_891; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_893 = 9'h176 == addrOdd[9:1] ? 32'h0 : _GEN_892; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_894 = 9'h177 == addrOdd[9:1] ? 32'h0 : _GEN_893; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_895 = 9'h178 == addrOdd[9:1] ? 32'h0 : _GEN_894; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_896 = 9'h179 == addrOdd[9:1] ? 32'h0 : _GEN_895; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_897 = 9'h17a == addrOdd[9:1] ? 32'h0 : _GEN_896; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_898 = 9'h17b == addrOdd[9:1] ? 32'h0 : _GEN_897; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_899 = 9'h17c == addrOdd[9:1] ? 32'h0 : _GEN_898; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_900 = 9'h17d == addrOdd[9:1] ? 32'h0 : _GEN_899; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_901 = 9'h17e == addrOdd[9:1] ? 32'h0 : _GEN_900; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_902 = 9'h17f == addrOdd[9:1] ? 32'h0 : _GEN_901; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_903 = 9'h180 == addrOdd[9:1] ? 32'h0 : _GEN_902; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_904 = 9'h181 == addrOdd[9:1] ? 32'h0 : _GEN_903; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_905 = 9'h182 == addrOdd[9:1] ? 32'h0 : _GEN_904; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_906 = 9'h183 == addrOdd[9:1] ? 32'h0 : _GEN_905; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_907 = 9'h184 == addrOdd[9:1] ? 32'h0 : _GEN_906; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_908 = 9'h185 == addrOdd[9:1] ? 32'h0 : _GEN_907; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_909 = 9'h186 == addrOdd[9:1] ? 32'h0 : _GEN_908; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_910 = 9'h187 == addrOdd[9:1] ? 32'h0 : _GEN_909; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_911 = 9'h188 == addrOdd[9:1] ? 32'h0 : _GEN_910; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_912 = 9'h189 == addrOdd[9:1] ? 32'h0 : _GEN_911; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_913 = 9'h18a == addrOdd[9:1] ? 32'h0 : _GEN_912; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_914 = 9'h18b == addrOdd[9:1] ? 32'h0 : _GEN_913; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_915 = 9'h18c == addrOdd[9:1] ? 32'h0 : _GEN_914; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_916 = 9'h18d == addrOdd[9:1] ? 32'h0 : _GEN_915; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_917 = 9'h18e == addrOdd[9:1] ? 32'h0 : _GEN_916; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_918 = 9'h18f == addrOdd[9:1] ? 32'h0 : _GEN_917; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_919 = 9'h190 == addrOdd[9:1] ? 32'h0 : _GEN_918; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_920 = 9'h191 == addrOdd[9:1] ? 32'h0 : _GEN_919; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_921 = 9'h192 == addrOdd[9:1] ? 32'h0 : _GEN_920; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_922 = 9'h193 == addrOdd[9:1] ? 32'h0 : _GEN_921; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_923 = 9'h194 == addrOdd[9:1] ? 32'h0 : _GEN_922; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_924 = 9'h195 == addrOdd[9:1] ? 32'h0 : _GEN_923; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_925 = 9'h196 == addrOdd[9:1] ? 32'h0 : _GEN_924; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_926 = 9'h197 == addrOdd[9:1] ? 32'h0 : _GEN_925; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_927 = 9'h198 == addrOdd[9:1] ? 32'h0 : _GEN_926; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_928 = 9'h199 == addrOdd[9:1] ? 32'h0 : _GEN_927; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_929 = 9'h19a == addrOdd[9:1] ? 32'h0 : _GEN_928; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_930 = 9'h19b == addrOdd[9:1] ? 32'h0 : _GEN_929; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_931 = 9'h19c == addrOdd[9:1] ? 32'h0 : _GEN_930; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_932 = 9'h19d == addrOdd[9:1] ? 32'h0 : _GEN_931; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_933 = 9'h19e == addrOdd[9:1] ? 32'h0 : _GEN_932; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_934 = 9'h19f == addrOdd[9:1] ? 32'h0 : _GEN_933; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_935 = 9'h1a0 == addrOdd[9:1] ? 32'h0 : _GEN_934; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_936 = 9'h1a1 == addrOdd[9:1] ? 32'h0 : _GEN_935; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_937 = 9'h1a2 == addrOdd[9:1] ? 32'h0 : _GEN_936; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_938 = 9'h1a3 == addrOdd[9:1] ? 32'h0 : _GEN_937; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_939 = 9'h1a4 == addrOdd[9:1] ? 32'h0 : _GEN_938; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_940 = 9'h1a5 == addrOdd[9:1] ? 32'h0 : _GEN_939; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_941 = 9'h1a6 == addrOdd[9:1] ? 32'h0 : _GEN_940; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_942 = 9'h1a7 == addrOdd[9:1] ? 32'h0 : _GEN_941; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_943 = 9'h1a8 == addrOdd[9:1] ? 32'h0 : _GEN_942; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_944 = 9'h1a9 == addrOdd[9:1] ? 32'h0 : _GEN_943; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_945 = 9'h1aa == addrOdd[9:1] ? 32'h0 : _GEN_944; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_946 = 9'h1ab == addrOdd[9:1] ? 32'h0 : _GEN_945; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_947 = 9'h1ac == addrOdd[9:1] ? 32'h0 : _GEN_946; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_948 = 9'h1ad == addrOdd[9:1] ? 32'h0 : _GEN_947; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_949 = 9'h1ae == addrOdd[9:1] ? 32'h0 : _GEN_948; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_950 = 9'h1af == addrOdd[9:1] ? 32'h0 : _GEN_949; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_951 = 9'h1b0 == addrOdd[9:1] ? 32'h0 : _GEN_950; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_952 = 9'h1b1 == addrOdd[9:1] ? 32'h0 : _GEN_951; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_953 = 9'h1b2 == addrOdd[9:1] ? 32'h0 : _GEN_952; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_954 = 9'h1b3 == addrOdd[9:1] ? 32'h0 : _GEN_953; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_955 = 9'h1b4 == addrOdd[9:1] ? 32'h0 : _GEN_954; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_956 = 9'h1b5 == addrOdd[9:1] ? 32'h0 : _GEN_955; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_957 = 9'h1b6 == addrOdd[9:1] ? 32'h0 : _GEN_956; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_958 = 9'h1b7 == addrOdd[9:1] ? 32'h0 : _GEN_957; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_959 = 9'h1b8 == addrOdd[9:1] ? 32'h0 : _GEN_958; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_960 = 9'h1b9 == addrOdd[9:1] ? 32'h0 : _GEN_959; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_961 = 9'h1ba == addrOdd[9:1] ? 32'h0 : _GEN_960; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_962 = 9'h1bb == addrOdd[9:1] ? 32'h0 : _GEN_961; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_963 = 9'h1bc == addrOdd[9:1] ? 32'h0 : _GEN_962; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_964 = 9'h1bd == addrOdd[9:1] ? 32'h0 : _GEN_963; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_965 = 9'h1be == addrOdd[9:1] ? 32'h0 : _GEN_964; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_966 = 9'h1bf == addrOdd[9:1] ? 32'h0 : _GEN_965; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_967 = 9'h1c0 == addrOdd[9:1] ? 32'h0 : _GEN_966; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_968 = 9'h1c1 == addrOdd[9:1] ? 32'h0 : _GEN_967; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_969 = 9'h1c2 == addrOdd[9:1] ? 32'h0 : _GEN_968; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_970 = 9'h1c3 == addrOdd[9:1] ? 32'h0 : _GEN_969; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_971 = 9'h1c4 == addrOdd[9:1] ? 32'h0 : _GEN_970; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_972 = 9'h1c5 == addrOdd[9:1] ? 32'h0 : _GEN_971; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_973 = 9'h1c6 == addrOdd[9:1] ? 32'h0 : _GEN_972; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_974 = 9'h1c7 == addrOdd[9:1] ? 32'h0 : _GEN_973; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_975 = 9'h1c8 == addrOdd[9:1] ? 32'h0 : _GEN_974; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_976 = 9'h1c9 == addrOdd[9:1] ? 32'h0 : _GEN_975; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_977 = 9'h1ca == addrOdd[9:1] ? 32'h0 : _GEN_976; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_978 = 9'h1cb == addrOdd[9:1] ? 32'h0 : _GEN_977; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_979 = 9'h1cc == addrOdd[9:1] ? 32'h0 : _GEN_978; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_980 = 9'h1cd == addrOdd[9:1] ? 32'h0 : _GEN_979; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_981 = 9'h1ce == addrOdd[9:1] ? 32'h0 : _GEN_980; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_982 = 9'h1cf == addrOdd[9:1] ? 32'h0 : _GEN_981; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_983 = 9'h1d0 == addrOdd[9:1] ? 32'h0 : _GEN_982; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_984 = 9'h1d1 == addrOdd[9:1] ? 32'h0 : _GEN_983; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_985 = 9'h1d2 == addrOdd[9:1] ? 32'h0 : _GEN_984; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_986 = 9'h1d3 == addrOdd[9:1] ? 32'h0 : _GEN_985; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_987 = 9'h1d4 == addrOdd[9:1] ? 32'h0 : _GEN_986; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_988 = 9'h1d5 == addrOdd[9:1] ? 32'h0 : _GEN_987; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_989 = 9'h1d6 == addrOdd[9:1] ? 32'h0 : _GEN_988; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_990 = 9'h1d7 == addrOdd[9:1] ? 32'h0 : _GEN_989; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_991 = 9'h1d8 == addrOdd[9:1] ? 32'h0 : _GEN_990; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_992 = 9'h1d9 == addrOdd[9:1] ? 32'h0 : _GEN_991; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_993 = 9'h1da == addrOdd[9:1] ? 32'h0 : _GEN_992; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_994 = 9'h1db == addrOdd[9:1] ? 32'h0 : _GEN_993; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_995 = 9'h1dc == addrOdd[9:1] ? 32'h0 : _GEN_994; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_996 = 9'h1dd == addrOdd[9:1] ? 32'h0 : _GEN_995; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_997 = 9'h1de == addrOdd[9:1] ? 32'h0 : _GEN_996; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_998 = 9'h1df == addrOdd[9:1] ? 32'h0 : _GEN_997; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_999 = 9'h1e0 == addrOdd[9:1] ? 32'h0 : _GEN_998; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1000 = 9'h1e1 == addrOdd[9:1] ? 32'h0 : _GEN_999; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1001 = 9'h1e2 == addrOdd[9:1] ? 32'h0 : _GEN_1000; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1002 = 9'h1e3 == addrOdd[9:1] ? 32'h0 : _GEN_1001; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1003 = 9'h1e4 == addrOdd[9:1] ? 32'h0 : _GEN_1002; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1004 = 9'h1e5 == addrOdd[9:1] ? 32'h0 : _GEN_1003; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1005 = 9'h1e6 == addrOdd[9:1] ? 32'h0 : _GEN_1004; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1006 = 9'h1e7 == addrOdd[9:1] ? 32'h0 : _GEN_1005; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1007 = 9'h1e8 == addrOdd[9:1] ? 32'h0 : _GEN_1006; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1008 = 9'h1e9 == addrOdd[9:1] ? 32'h0 : _GEN_1007; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1009 = 9'h1ea == addrOdd[9:1] ? 32'h0 : _GEN_1008; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1010 = 9'h1eb == addrOdd[9:1] ? 32'h0 : _GEN_1009; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1011 = 9'h1ec == addrOdd[9:1] ? 32'h0 : _GEN_1010; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1012 = 9'h1ed == addrOdd[9:1] ? 32'h0 : _GEN_1011; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1013 = 9'h1ee == addrOdd[9:1] ? 32'h0 : _GEN_1012; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1014 = 9'h1ef == addrOdd[9:1] ? 32'h0 : _GEN_1013; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1015 = 9'h1f0 == addrOdd[9:1] ? 32'h0 : _GEN_1014; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1016 = 9'h1f1 == addrOdd[9:1] ? 32'h0 : _GEN_1015; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1017 = 9'h1f2 == addrOdd[9:1] ? 32'h0 : _GEN_1016; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1018 = 9'h1f3 == addrOdd[9:1] ? 32'h0 : _GEN_1017; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1019 = 9'h1f4 == addrOdd[9:1] ? 32'h0 : _GEN_1018; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1020 = 9'h1f5 == addrOdd[9:1] ? 32'h0 : _GEN_1019; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1021 = 9'h1f6 == addrOdd[9:1] ? 32'h0 : _GEN_1020; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1022 = 9'h1f7 == addrOdd[9:1] ? 32'h0 : _GEN_1021; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1023 = 9'h1f8 == addrOdd[9:1] ? 32'h0 : _GEN_1022; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1024 = 9'h1f9 == addrOdd[9:1] ? 32'h0 : _GEN_1023; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1025 = 9'h1fa == addrOdd[9:1] ? 32'h0 : _GEN_1024; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] _GEN_1026 = 9'h1fb == addrOdd[9:1] ? 32'h0 : _GEN_1025; // @[Fetch.scala 101:25 Fetch.scala 101:25]
  wire [31:0] instr_b_rom = _T_14 ? data_odd : data_even; // @[Fetch.scala 103:24]
  wire [31:0] instr_b_cache = _T_14 ? io_icachefe_instrOdd : io_icachefe_instrEven; // @[Fetch.scala 107:26]
  wire [31:0] _T_32 = selCache ? instr_b_cache : instr_b_rom; // @[Fetch.scala 113:24]
  wire [29:0] pcNext = pc_next; // @[Fetch.scala 119:8]
  wire [29:0] _GEN_1034 = {{19'd0}, relBaseReg}; // @[Fetch.scala 138:21]
  wire [29:0] relPc = pcReg - _GEN_1034; // @[Fetch.scala 138:21]
  wire [29:0] _T_56 = relPc + 30'h2; // @[Fetch.scala 147:36]
  wire [29:0] _T_58 = relPc + 30'h1; // @[Fetch.scala 147:53]
  wire  selSpmNext = io_ena ? io_icachefe_memSel[1] : selSpm; // @[Fetch.scala 73:17 Fetch.scala 74:16 Fetch.scala 69:14]
  wire  selCacheNext = io_ena ? io_icachefe_memSel[0] : selCache; // @[Fetch.scala 73:17 Fetch.scala 75:18 Fetch.scala 71:16]
  wire [10:0] relBaseNext = io_ena ? _GEN_2 : relBaseReg; // @[Fetch.scala 89:16 Fetch.scala 85:15]
  wire [31:0] relocNext = io_ena ? _GEN_3 : relocReg; // @[Fetch.scala 89:16 Fetch.scala 87:13]
  MemBlock_2 MemBlock ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_clock),
    .io_rdAddr(MemBlock_io_rdAddr),
    .io_rdData(MemBlock_io_rdData),
    .io_wrAddr(MemBlock_io_wrAddr),
    .io_wrEna(MemBlock_io_wrEna),
    .io_wrData(MemBlock_io_wrData)
  );
  MemBlock_2 MemBlock_1 ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_1_clock),
    .io_rdAddr(MemBlock_1_io_rdAddr),
    .io_rdData(MemBlock_1_io_rdData),
    .io_wrAddr(MemBlock_1_io_wrAddr),
    .io_wrEna(MemBlock_1_io_wrEna),
    .io_wrData(MemBlock_1_io_wrData)
  );
  assign io_fedec_instr_a = selSpm ? instr_a_ispm : _T_31; // @[Fetch.scala 110:20]
  assign io_fedec_instr_b = selSpm ? instr_b_ispm : _T_32; // @[Fetch.scala 112:20]
  assign io_fedec_pc = pcReg; // @[Fetch.scala 140:15]
  assign io_fedec_base = baseReg[29:0]; // @[Fetch.scala 141:17]
  assign io_fedec_reloc = relocReg; // @[Fetch.scala 142:18]
  assign io_fedec_relPc = pcReg - _GEN_1034; // @[Fetch.scala 138:21]
  assign io_feex_pc = b_valid ? _T_56 : _T_58; // @[Fetch.scala 147:20]
  assign io_feicache_addrEven = {{2'd0}, addrEven}; // @[Fetch.scala 132:26 Fetch.scala 133:14 Fetch.scala 130:12]
  assign io_feicache_addrOdd = {{2'd0}, addrOdd}; // @[Fetch.scala 132:26 Fetch.scala 134:13 Fetch.scala 131:11]
  assign MemBlock_clock = clock;
  assign MemBlock_io_rdAddr = addrEven[7:1]; // @[Fetch.scala 55:40]
  assign MemBlock_io_wrAddr = io_memfe_addr[9:3]; // @[Fetch.scala 51:41]
  assign MemBlock_io_wrEna = _T_2 & ~io_memfe_addr[2]; // @[Fetch.scala 49:27]
  assign MemBlock_io_wrData = io_memfe_data; // @[MemBlock.scala 36:12]
  assign MemBlock_1_clock = clock;
  assign MemBlock_1_io_rdAddr = addrOdd[7:1]; // @[Fetch.scala 56:37]
  assign MemBlock_1_io_wrAddr = io_memfe_addr[9:3]; // @[Fetch.scala 52:39]
  assign MemBlock_1_io_wrEna = _T_2 & io_memfe_addr[2]; // @[Fetch.scala 50:26]
  assign MemBlock_1_io_wrData = io_memfe_data; // @[MemBlock.scala 36:12]
  always @(posedge clock) begin
    if (reset) begin // @[Fetch.scala 21:22]
      pcReg <= 30'h1; // @[Fetch.scala 21:22]
    end else if (io_ena & ~reset) begin // @[Fetch.scala 132:26]
      pcReg <= pcNext; // @[Fetch.scala 135:11]
    end
    if (reset) begin // @[Fetch.scala 25:24]
      addrEvenReg <= 30'h2; // @[Fetch.scala 25:24]
    end else if (io_ena & ~reset) begin // @[Fetch.scala 132:26]
      addrEvenReg <= _T_52; // @[Fetch.scala 133:14]
    end
    if (reset) begin // @[Fetch.scala 26:23]
      addrOddReg <= 30'h1; // @[Fetch.scala 26:23]
    end else if (io_ena & ~reset) begin // @[Fetch.scala 132:26]
      addrOddReg <= _T_53; // @[Fetch.scala 134:13]
    end
    if (reset) begin // @[Fetch.scala 65:23]
      selSpm <= 1'h0; // @[Fetch.scala 65:23]
    end else if (io_ena) begin // @[Fetch.scala 73:17]
      selSpm <= io_icachefe_memSel[1]; // @[Fetch.scala 74:16]
    end
    if (reset) begin // @[Fetch.scala 66:25]
      selCache <= 1'h0; // @[Fetch.scala 66:25]
    end else if (io_ena) begin // @[Fetch.scala 73:17]
      selCache <= io_icachefe_memSel[0]; // @[Fetch.scala 75:18]
    end
    if (9'h1ff == addrEven[9:1]) begin // @[Fetch.scala 100:26]
      data_even <= 32'h0; // @[Fetch.scala 100:26]
    end else if (9'h1fe == addrEven[9:1]) begin // @[Fetch.scala 100:26]
      data_even <= 32'h0; // @[Fetch.scala 100:26]
    end else if (9'h1fd == addrEven[9:1]) begin // @[Fetch.scala 100:26]
      data_even <= 32'h0; // @[Fetch.scala 100:26]
    end else if (9'h1fc == addrEven[9:1]) begin // @[Fetch.scala 100:26]
      data_even <= 32'h0; // @[Fetch.scala 100:26]
    end else begin
      data_even <= _GEN_514;
    end
    if (9'h1ff == addrOdd[9:1]) begin // @[Fetch.scala 101:25]
      data_odd <= 32'h0; // @[Fetch.scala 101:25]
    end else if (9'h1fe == addrOdd[9:1]) begin // @[Fetch.scala 101:25]
      data_odd <= 32'h0; // @[Fetch.scala 101:25]
    end else if (9'h1fd == addrOdd[9:1]) begin // @[Fetch.scala 101:25]
      data_odd <= 32'h0; // @[Fetch.scala 101:25]
    end else if (9'h1fc == addrOdd[9:1]) begin // @[Fetch.scala 101:25]
      data_odd <= 32'h0; // @[Fetch.scala 101:25]
    end else begin
      data_odd <= _GEN_1026;
    end
    if (reset) begin // @[Fetch.scala 79:24]
      baseReg <= 32'h0; // @[Fetch.scala 79:24]
    end else if (io_ena) begin // @[Fetch.scala 89:16]
      baseReg <= io_icachefe_base; // @[Fetch.scala 90:13]
    end
    if (reset) begin // @[Fetch.scala 80:27]
      relBaseReg <= 11'h1; // @[Fetch.scala 80:27]
    end else if (io_ena) begin // @[Fetch.scala 89:16]
      if (io_memfe_doCallRet) begin // @[Fetch.scala 91:31]
        relBaseReg <= io_icachefe_relBase; // @[Fetch.scala 92:19]
      end
    end
    if (reset) begin // @[Fetch.scala 81:25]
      relocReg <= 32'h0; // @[Fetch.scala 81:25]
    end else if (io_ena) begin // @[Fetch.scala 89:16]
      if (io_memfe_doCallRet) begin // @[Fetch.scala 91:31]
        relocReg <= io_icachefe_reloc; // @[Fetch.scala 93:17]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pcReg = _RAND_0[29:0];
  _RAND_1 = {1{`RANDOM}};
  addrEvenReg = _RAND_1[29:0];
  _RAND_2 = {1{`RANDOM}};
  addrOddReg = _RAND_2[29:0];
  _RAND_3 = {1{`RANDOM}};
  selSpm = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  selCache = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  data_even = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  data_odd = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  baseReg = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  relBaseReg = _RAND_8[10:0];
  _RAND_9 = {1{`RANDOM}};
  relocReg = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegisterFile(
  input         clock,
  input         io_ena,
  input  [4:0]  io_rfRead_rsAddr_0,
  input  [4:0]  io_rfRead_rsAddr_1,
  input  [4:0]  io_rfRead_rsAddr_2,
  input  [4:0]  io_rfRead_rsAddr_3,
  output [31:0] io_rfRead_rsData_0,
  output [31:0] io_rfRead_rsData_1,
  output [31:0] io_rfRead_rsData_2,
  output [31:0] io_rfRead_rsData_3,
  input  [4:0]  io_rfWrite_0_addr,
  input  [31:0] io_rfWrite_0_data,
  input         io_rfWrite_0_valid,
  input  [4:0]  io_rfWrite_1_addr,
  input  [31:0] io_rfWrite_1_data,
  input         io_rfWrite_1_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] rf [0:31];
  wire [31:0] rf_MPORT_data;
  wire [4:0] rf_MPORT_addr;
  wire [31:0] rf_MPORT_1_data;
  wire [4:0] rf_MPORT_1_addr;
  wire [31:0] rf_MPORT_2_data;
  wire [4:0] rf_MPORT_2_addr;
  wire [31:0] rf_MPORT_3_data;
  wire [4:0] rf_MPORT_3_addr;
  wire [31:0] rf_MPORT_4_data;
  wire [4:0] rf_MPORT_4_addr;
  wire  rf_MPORT_4_mask;
  wire  rf_MPORT_4_en;
  wire [31:0] rf_MPORT_5_data;
  wire [4:0] rf_MPORT_5_addr;
  wire  rf_MPORT_5_mask;
  wire  rf_MPORT_5_en;
  reg [4:0] addrReg_0; // @[RegisterFile.scala 22:20]
  reg [4:0] addrReg_1; // @[RegisterFile.scala 22:20]
  reg [4:0] addrReg_2; // @[RegisterFile.scala 22:20]
  reg [4:0] addrReg_3; // @[RegisterFile.scala 22:20]
  reg [31:0] wrReg_0_data; // @[RegisterFile.scala 23:20]
  reg [31:0] wrReg_1_data; // @[RegisterFile.scala 23:20]
  reg  fwReg_0_0; // @[RegisterFile.scala 24:20]
  reg  fwReg_0_1; // @[RegisterFile.scala 24:20]
  reg  fwReg_1_0; // @[RegisterFile.scala 24:20]
  reg  fwReg_1_1; // @[RegisterFile.scala 24:20]
  reg  fwReg_2_0; // @[RegisterFile.scala 24:20]
  reg  fwReg_2_1; // @[RegisterFile.scala 24:20]
  reg  fwReg_3_0; // @[RegisterFile.scala 24:20]
  reg  fwReg_3_1; // @[RegisterFile.scala 24:20]
  wire [31:0] _GEN_18 = fwReg_0_0 ? wrReg_0_data : rf_MPORT_data; // @[RegisterFile.scala 40:26 RegisterFile.scala 41:29 RegisterFile.scala 38:25]
  wire [31:0] _GEN_19 = fwReg_0_1 ? wrReg_1_data : _GEN_18; // @[RegisterFile.scala 40:26 RegisterFile.scala 41:29]
  wire [31:0] _GEN_21 = fwReg_1_0 ? wrReg_0_data : rf_MPORT_1_data; // @[RegisterFile.scala 40:26 RegisterFile.scala 41:29 RegisterFile.scala 38:25]
  wire [31:0] _GEN_22 = fwReg_1_1 ? wrReg_1_data : _GEN_21; // @[RegisterFile.scala 40:26 RegisterFile.scala 41:29]
  wire [31:0] _GEN_24 = fwReg_2_0 ? wrReg_0_data : rf_MPORT_2_data; // @[RegisterFile.scala 40:26 RegisterFile.scala 41:29 RegisterFile.scala 38:25]
  wire [31:0] _GEN_25 = fwReg_2_1 ? wrReg_1_data : _GEN_24; // @[RegisterFile.scala 40:26 RegisterFile.scala 41:29]
  wire [31:0] _GEN_27 = fwReg_3_0 ? wrReg_0_data : rf_MPORT_3_data; // @[RegisterFile.scala 40:26 RegisterFile.scala 41:29 RegisterFile.scala 38:25]
  wire [31:0] _GEN_28 = fwReg_3_1 ? wrReg_1_data : _GEN_27; // @[RegisterFile.scala 40:26 RegisterFile.scala 41:29]
  assign rf_MPORT_addr = addrReg_0;
  assign rf_MPORT_data = rf[rf_MPORT_addr];
  assign rf_MPORT_1_addr = addrReg_1;
  assign rf_MPORT_1_data = rf[rf_MPORT_1_addr];
  assign rf_MPORT_2_addr = addrReg_2;
  assign rf_MPORT_2_data = rf[rf_MPORT_2_addr];
  assign rf_MPORT_3_addr = addrReg_3;
  assign rf_MPORT_3_data = rf[rf_MPORT_3_addr];
  assign rf_MPORT_4_data = io_rfWrite_1_data;
  assign rf_MPORT_4_addr = io_rfWrite_1_addr;
  assign rf_MPORT_4_mask = 1'h1;
  assign rf_MPORT_4_en = io_rfWrite_1_valid;
  assign rf_MPORT_5_data = io_rfWrite_0_data;
  assign rf_MPORT_5_addr = io_rfWrite_0_addr;
  assign rf_MPORT_5_mask = 1'h1;
  assign rf_MPORT_5_en = io_rfWrite_0_valid;
  assign io_rfRead_rsData_0 = addrReg_0 == 5'h0 ? 32'h0 : _GEN_19; // @[RegisterFile.scala 44:34 RegisterFile.scala 45:27]
  assign io_rfRead_rsData_1 = addrReg_1 == 5'h0 ? 32'h0 : _GEN_22; // @[RegisterFile.scala 44:34 RegisterFile.scala 45:27]
  assign io_rfRead_rsData_2 = addrReg_2 == 5'h0 ? 32'h0 : _GEN_25; // @[RegisterFile.scala 44:34 RegisterFile.scala 45:27]
  assign io_rfRead_rsData_3 = addrReg_3 == 5'h0 ? 32'h0 : _GEN_28; // @[RegisterFile.scala 44:34 RegisterFile.scala 45:27]
  always @(posedge clock) begin
    if(rf_MPORT_4_en & rf_MPORT_4_mask) begin
      rf[rf_MPORT_4_addr] <= rf_MPORT_4_data;
    end
    if(rf_MPORT_5_en & rf_MPORT_5_mask) begin
      rf[rf_MPORT_5_addr] <= rf_MPORT_5_data;
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      addrReg_0 <= io_rfRead_rsAddr_0; // @[RegisterFile.scala 27:13]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      addrReg_1 <= io_rfRead_rsAddr_1; // @[RegisterFile.scala 27:13]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      addrReg_2 <= io_rfRead_rsAddr_2; // @[RegisterFile.scala 27:13]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      addrReg_3 <= io_rfRead_rsAddr_3; // @[RegisterFile.scala 27:13]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      wrReg_0_data <= io_rfWrite_0_data; // @[RegisterFile.scala 28:11]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      wrReg_1_data <= io_rfWrite_1_data; // @[RegisterFile.scala 28:11]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      fwReg_0_0 <= io_rfRead_rsAddr_0 == io_rfWrite_0_addr & io_rfWrite_0_valid; // @[RegisterFile.scala 31:21]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      fwReg_0_1 <= io_rfRead_rsAddr_0 == io_rfWrite_1_addr & io_rfWrite_1_valid; // @[RegisterFile.scala 31:21]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      fwReg_1_0 <= io_rfRead_rsAddr_1 == io_rfWrite_0_addr & io_rfWrite_0_valid; // @[RegisterFile.scala 31:21]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      fwReg_1_1 <= io_rfRead_rsAddr_1 == io_rfWrite_1_addr & io_rfWrite_1_valid; // @[RegisterFile.scala 31:21]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      fwReg_2_0 <= io_rfRead_rsAddr_2 == io_rfWrite_0_addr & io_rfWrite_0_valid; // @[RegisterFile.scala 31:21]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      fwReg_2_1 <= io_rfRead_rsAddr_2 == io_rfWrite_1_addr & io_rfWrite_1_valid; // @[RegisterFile.scala 31:21]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      fwReg_3_0 <= io_rfRead_rsAddr_3 == io_rfWrite_0_addr & io_rfWrite_0_valid; // @[RegisterFile.scala 31:21]
    end
    if (io_ena) begin // @[RegisterFile.scala 26:17]
      fwReg_3_1 <= io_rfRead_rsAddr_3 == io_rfWrite_1_addr & io_rfWrite_1_valid; // @[RegisterFile.scala 31:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    rf[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  addrReg_0 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  addrReg_1 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  addrReg_2 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  addrReg_3 = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  wrReg_0_data = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  wrReg_1_data = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  fwReg_0_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  fwReg_0_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  fwReg_1_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  fwReg_1_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  fwReg_2_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  fwReg_2_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  fwReg_3_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  fwReg_3_1 = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decode(
  input         clock,
  input         reset,
  input         io_ena,
  input         io_flush,
  input  [31:0] io_fedec_instr_a,
  input  [31:0] io_fedec_instr_b,
  input  [29:0] io_fedec_pc,
  input  [29:0] io_fedec_base,
  input  [31:0] io_fedec_reloc,
  input  [29:0] io_fedec_relPc,
  output [29:0] io_decex_base,
  output [29:0] io_decex_relPc,
  output [3:0]  io_decex_pred_0,
  output [3:0]  io_decex_pred_1,
  output [3:0]  io_decex_aluOp_0_func,
  output        io_decex_aluOp_0_isMul,
  output        io_decex_aluOp_0_isCmp,
  output        io_decex_aluOp_0_isPred,
  output        io_decex_aluOp_0_isBCpy,
  output        io_decex_aluOp_0_isMTS,
  output        io_decex_aluOp_0_isMFS,
  output [3:0]  io_decex_aluOp_1_func,
  output        io_decex_aluOp_1_isCmp,
  output        io_decex_aluOp_1_isPred,
  output        io_decex_aluOp_1_isBCpy,
  output        io_decex_aluOp_1_isMTS,
  output        io_decex_aluOp_1_isMFS,
  output [1:0]  io_decex_predOp_0_func,
  output [2:0]  io_decex_predOp_0_dest,
  output [3:0]  io_decex_predOp_0_s1Addr,
  output [3:0]  io_decex_predOp_0_s2Addr,
  output [1:0]  io_decex_predOp_1_func,
  output [2:0]  io_decex_predOp_1_dest,
  output [3:0]  io_decex_predOp_1_s1Addr,
  output [3:0]  io_decex_predOp_1_s2Addr,
  output        io_decex_jmpOp_branch,
  output [29:0] io_decex_jmpOp_target,
  output [31:0] io_decex_jmpOp_reloc,
  output        io_decex_memOp_load,
  output        io_decex_memOp_store,
  output        io_decex_memOp_hword,
  output        io_decex_memOp_byte,
  output        io_decex_memOp_zext,
  output [1:0]  io_decex_memOp_typ,
  output [2:0]  io_decex_stackOp,
  output [4:0]  io_decex_rsAddr_0,
  output [4:0]  io_decex_rsAddr_1,
  output [4:0]  io_decex_rsAddr_2,
  output [4:0]  io_decex_rsAddr_3,
  output [31:0] io_decex_rsData_0,
  output [31:0] io_decex_rsData_1,
  output [31:0] io_decex_rsData_2,
  output [31:0] io_decex_rsData_3,
  output [4:0]  io_decex_rdAddr_0,
  output [4:0]  io_decex_rdAddr_1,
  output [31:0] io_decex_immVal_0,
  output [31:0] io_decex_immVal_1,
  output        io_decex_immOp_0,
  output        io_decex_immOp_1,
  output        io_decex_wrRd_0,
  output        io_decex_wrRd_1,
  output [31:0] io_decex_callAddr,
  output        io_decex_call,
  output        io_decex_ret,
  output        io_decex_brcf,
  output        io_decex_trap,
  output        io_decex_xcall,
  output        io_decex_xret,
  output [4:0]  io_decex_xsrc,
  output        io_decex_nonDelayed,
  output        io_decex_illOp,
  input  [4:0]  io_rfWrite_0_addr,
  input  [31:0] io_rfWrite_0_data,
  input         io_rfWrite_0_valid,
  input  [4:0]  io_rfWrite_1_addr,
  input  [31:0] io_rfWrite_1_data,
  input         io_rfWrite_1_valid,
  input         io_exc_exc,
  input  [29:0] io_exc_excBase,
  input  [29:0] io_exc_excAddr,
  input         io_exc_intr,
  input  [31:0] io_exc_addr,
  input  [4:0]  io_exc_src,
  input         io_exc_local
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  rf_clock; // @[Decode.scala 19:18]
  wire  rf_io_ena; // @[Decode.scala 19:18]
  wire [4:0] rf_io_rfRead_rsAddr_0; // @[Decode.scala 19:18]
  wire [4:0] rf_io_rfRead_rsAddr_1; // @[Decode.scala 19:18]
  wire [4:0] rf_io_rfRead_rsAddr_2; // @[Decode.scala 19:18]
  wire [4:0] rf_io_rfRead_rsAddr_3; // @[Decode.scala 19:18]
  wire [31:0] rf_io_rfRead_rsData_0; // @[Decode.scala 19:18]
  wire [31:0] rf_io_rfRead_rsData_1; // @[Decode.scala 19:18]
  wire [31:0] rf_io_rfRead_rsData_2; // @[Decode.scala 19:18]
  wire [31:0] rf_io_rfRead_rsData_3; // @[Decode.scala 19:18]
  wire [4:0] rf_io_rfWrite_0_addr; // @[Decode.scala 19:18]
  wire [31:0] rf_io_rfWrite_0_data; // @[Decode.scala 19:18]
  wire  rf_io_rfWrite_0_valid; // @[Decode.scala 19:18]
  wire [4:0] rf_io_rfWrite_1_addr; // @[Decode.scala 19:18]
  wire [31:0] rf_io_rfWrite_1_data; // @[Decode.scala 19:18]
  wire  rf_io_rfWrite_1_valid; // @[Decode.scala 19:18]
  reg [31:0] decReg_instr_a; // @[Decode.scala 32:19]
  reg [31:0] decReg_instr_b; // @[Decode.scala 32:19]
  reg [29:0] decReg_pc; // @[Decode.scala 32:19]
  reg [29:0] decReg_base; // @[Decode.scala 32:19]
  reg [31:0] decReg_reloc; // @[Decode.scala 32:19]
  reg [29:0] decReg_relPc; // @[Decode.scala 32:19]
  wire  dual = decReg_instr_a[31] & decReg_instr_a[26:22] != 5'h1f; // @[Decode.scala 63:46]
  wire [11:0] lo = decReg_instr_a[11:0]; // @[Decode.scala 72:33]
  wire [12:0] _T_15 = {1'h0,lo}; // @[Cat.scala 30:58]
  wire  _T_18 = decReg_instr_a[26:25] == 2'h0; // @[Decode.scala 78:23]
  wire [2:0] lo_1 = decReg_instr_a[24:22]; // @[Decode.scala 79:51]
  wire [3:0] _T_19 = {1'h0,lo_1}; // @[Cat.scala 30:58]
  wire [3:0] _GEN_9 = decReg_instr_a[26:25] == 2'h0 ? _T_19 : decReg_instr_a[3:0]; // @[Decode.scala 78:40 Decode.scala 79:30 Decode.scala 75:28]
  wire  _T_21 = 3'h0 == decReg_instr_a[6:4]; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h1 == decReg_instr_a[6:4]; // @[Conditional.scala 37:30]
  wire  _T_23 = 3'h2 == decReg_instr_a[6:4]; // @[Conditional.scala 37:30]
  wire  _T_24 = 3'h3 == decReg_instr_a[6:4]; // @[Conditional.scala 37:30]
  wire  _T_25 = 3'h6 == decReg_instr_a[6:4]; // @[Conditional.scala 37:30]
  wire [5:0] _T_26 = {1'h0,decReg_instr_a[11:7]}; // @[Cat.scala 30:58]
  wire  _T_27 = 3'h4 == decReg_instr_a[6:4]; // @[Conditional.scala 37:30]
  wire  _T_28 = 3'h5 == decReg_instr_a[6:4]; // @[Conditional.scala 37:30]
  wire  _GEN_13 = _T_28 | _T_18; // @[Conditional.scala 39:67 Decode.scala 114:28]
  wire [12:0] _GEN_16 = _T_28 ? {{7'd0}, _T_26} : _T_15; // @[Conditional.scala 39:67 Decode.scala 117:18 Decode.scala 72:12]
  wire  _GEN_19 = _T_27 | _GEN_13; // @[Conditional.scala 39:67 Decode.scala 111:22]
  wire  _GEN_20 = _T_27 ? _T_18 : _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_21 = _T_27 ? 1'h0 : _T_28; // @[Conditional.scala 39:67 connections.scala 50:12]
  wire [12:0] _GEN_23 = _T_27 ? _T_15 : _GEN_16; // @[Conditional.scala 39:67 Decode.scala 72:12]
  wire  _GEN_25 = _T_25 | _GEN_20; // @[Conditional.scala 39:67 Decode.scala 105:29]
  wire [12:0] _GEN_26 = _T_25 ? {{7'd0}, _T_26} : _GEN_23; // @[Conditional.scala 39:67 Decode.scala 106:18]
  wire  _GEN_27 = _T_25 | _GEN_19; // @[Conditional.scala 39:67 Decode.scala 107:22]
  wire  _GEN_28 = _T_25 ? 1'h0 : _T_27; // @[Conditional.scala 39:67 connections.scala 49:12]
  wire  _GEN_29 = _T_25 ? _T_18 : _GEN_20; // @[Conditional.scala 39:67]
  wire  _GEN_30 = _T_25 ? 1'h0 : _GEN_21; // @[Conditional.scala 39:67 connections.scala 50:12]
  wire  _GEN_31 = _T_24 | _T_25; // @[Conditional.scala 39:67 Decode.scala 100:35]
  wire  _GEN_32 = _T_24 | _GEN_27; // @[Conditional.scala 39:67 Decode.scala 101:22]
  wire  _GEN_33 = _T_24 ? _T_18 : _GEN_25; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_34 = _T_24 ? _T_15 : _GEN_26; // @[Conditional.scala 39:67 Decode.scala 72:12]
  wire  _GEN_35 = _T_24 ? 1'h0 : _GEN_28; // @[Conditional.scala 39:67 connections.scala 49:12]
  wire  _GEN_36 = _T_24 ? _T_18 : _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_37 = _T_24 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67 connections.scala 50:12]
  wire  _GEN_39 = _T_23 | _GEN_32; // @[Conditional.scala 39:67 Decode.scala 97:22]
  wire  _GEN_40 = _T_23 ? 1'h0 : _GEN_31; // @[Conditional.scala 39:67 connections.scala 48:11]
  wire  _GEN_41 = _T_23 ? _T_18 : _GEN_33; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_42 = _T_23 ? _T_15 : _GEN_34; // @[Conditional.scala 39:67 Decode.scala 72:12]
  wire  _GEN_43 = _T_23 ? 1'h0 : _GEN_35; // @[Conditional.scala 39:67 connections.scala 49:12]
  wire  _GEN_44 = _T_23 ? _T_18 : _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_45 = _T_23 ? 1'h0 : _GEN_37; // @[Conditional.scala 39:67 connections.scala 50:12]
  wire  _GEN_46 = _T_22 | _GEN_44; // @[Conditional.scala 39:67 Decode.scala 92:28]
  wire  _GEN_47 = _T_22 | _GEN_39; // @[Conditional.scala 39:67 Decode.scala 93:22]
  wire  _GEN_48 = _T_22 ? 1'h0 : _T_23; // @[Conditional.scala 39:67 connections.scala 47:11]
  wire  _GEN_49 = _T_22 ? 1'h0 : _GEN_40; // @[Conditional.scala 39:67 connections.scala 48:11]
  wire  _GEN_50 = _T_22 ? _T_18 : _GEN_41; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_51 = _T_22 ? _T_15 : _GEN_42; // @[Conditional.scala 39:67 Decode.scala 72:12]
  wire  _GEN_52 = _T_22 ? 1'h0 : _GEN_43; // @[Conditional.scala 39:67 connections.scala 49:12]
  wire  _GEN_53 = _T_22 ? 1'h0 : _GEN_45; // @[Conditional.scala 39:67 connections.scala 50:12]
  wire  _GEN_54 = _T_21 | _GEN_46; // @[Conditional.scala 40:58 Decode.scala 88:28]
  wire  _GEN_55 = _T_21 | _GEN_47; // @[Conditional.scala 40:58 Decode.scala 89:22]
  wire  _GEN_56 = _T_21 ? 1'h0 : _GEN_48; // @[Conditional.scala 40:58 connections.scala 47:11]
  wire  _GEN_57 = _T_21 ? 1'h0 : _GEN_49; // @[Conditional.scala 40:58 connections.scala 48:11]
  wire  _GEN_58 = _T_21 ? _T_18 : _GEN_50; // @[Conditional.scala 40:58]
  wire [12:0] _GEN_59 = _T_21 ? _T_15 : _GEN_51; // @[Conditional.scala 40:58 Decode.scala 72:12]
  wire  _GEN_60 = _T_21 ? 1'h0 : _GEN_52; // @[Conditional.scala 40:58 connections.scala 49:12]
  wire  _GEN_61 = _T_21 ? 1'h0 : _GEN_53; // @[Conditional.scala 40:58 connections.scala 50:12]
  wire  _GEN_62 = decReg_instr_a[26:22] == 5'h8 ? _GEN_54 : _T_18; // @[Decode.scala 85:33]
  wire  _GEN_63 = decReg_instr_a[26:22] == 5'h8 ? _GEN_55 : _T_18; // @[Decode.scala 85:33]
  wire  _GEN_64 = decReg_instr_a[26:22] == 5'h8 & _GEN_56; // @[Decode.scala 85:33 connections.scala 47:11]
  wire  _GEN_65 = decReg_instr_a[26:22] == 5'h8 & _GEN_57; // @[Decode.scala 85:33 connections.scala 48:11]
  wire  _GEN_66 = decReg_instr_a[26:22] == 5'h8 ? _GEN_58 : _T_18; // @[Decode.scala 85:33]
  wire [12:0] _GEN_67 = decReg_instr_a[26:22] == 5'h8 ? _GEN_59 : _T_15; // @[Decode.scala 85:33 Decode.scala 72:12]
  wire  _GEN_68 = decReg_instr_a[26:22] == 5'h8 & _GEN_60; // @[Decode.scala 85:33 connections.scala 49:12]
  wire  _GEN_69 = decReg_instr_a[26:22] == 5'h8 & _GEN_61; // @[Decode.scala 85:33 connections.scala 50:12]
  wire  _GEN_71 = _T_24 | _GEN_62; // @[Conditional.scala 39:67 Decode.scala 131:28]
  wire  _GEN_72 = _T_24 | _GEN_63; // @[Conditional.scala 39:67 Decode.scala 132:22]
  wire  _GEN_74 = _T_23 | _GEN_72; // @[Conditional.scala 40:58 Decode.scala 127:22]
  wire  _GEN_75 = _T_23 ? 1'h0 : _T_24; // @[Conditional.scala 40:58 connections.scala 52:11]
  wire  _GEN_76 = _T_23 ? _GEN_62 : _GEN_71; // @[Conditional.scala 40:58]
  wire  _GEN_77 = decReg_instr_a[26:22] == 5'h9 & _T_23; // @[Decode.scala 123:33 connections.scala 51:11]
  wire  _GEN_78 = decReg_instr_a[26:22] == 5'h9 ? _GEN_74 : _GEN_63; // @[Decode.scala 123:33]
  wire  _GEN_79 = decReg_instr_a[26:22] == 5'h9 & _GEN_75; // @[Decode.scala 123:33 connections.scala 52:11]
  wire  _GEN_80 = decReg_instr_a[26:22] == 5'h9 ? _GEN_76 : _GEN_62; // @[Decode.scala 123:33]
  wire  hi = decReg_instr_a[3]; // @[Decode.scala 141:41]
  wire  lo_4 = decReg_instr_a[0]; // @[Decode.scala 141:51]
  wire [1:0] _T_33 = {hi,lo_4}; // @[Cat.scala 30:58]
  wire [11:0] lo_5 = decReg_instr_b[11:0]; // @[Decode.scala 72:33]
  wire [12:0] _T_41 = {1'h0,lo_5}; // @[Cat.scala 30:58]
  wire  _T_44 = decReg_instr_b[26:25] == 2'h0; // @[Decode.scala 78:23]
  wire [2:0] lo_6 = decReg_instr_b[24:22]; // @[Decode.scala 79:51]
  wire [3:0] _T_45 = {1'h0,lo_6}; // @[Cat.scala 30:58]
  wire [3:0] _GEN_81 = decReg_instr_b[26:25] == 2'h0 ? _T_45 : decReg_instr_b[3:0]; // @[Decode.scala 78:40 Decode.scala 79:30 Decode.scala 75:28]
  wire  _GEN_82 = decReg_instr_b[26:25] == 2'h0 & dual; // @[Decode.scala 78:40 Decode.scala 80:25 connections.scala 151:11]
  wire  _T_47 = 3'h0 == decReg_instr_b[6:4]; // @[Conditional.scala 37:30]
  wire  _T_48 = 3'h1 == decReg_instr_b[6:4]; // @[Conditional.scala 37:30]
  wire  _T_49 = 3'h2 == decReg_instr_b[6:4]; // @[Conditional.scala 37:30]
  wire  _T_50 = 3'h3 == decReg_instr_b[6:4]; // @[Conditional.scala 37:30]
  wire  _T_51 = 3'h6 == decReg_instr_b[6:4]; // @[Conditional.scala 37:30]
  wire [5:0] _T_52 = {1'h0,decReg_instr_b[11:7]}; // @[Cat.scala 30:58]
  wire  _T_53 = 3'h4 == decReg_instr_b[6:4]; // @[Conditional.scala 37:30]
  wire  _T_54 = 3'h5 == decReg_instr_b[6:4]; // @[Conditional.scala 37:30]
  wire  _GEN_85 = _T_54 ? dual : _GEN_82; // @[Conditional.scala 39:67 Decode.scala 114:28]
  wire  _GEN_86 = _T_54 & dual; // @[Conditional.scala 39:67 Decode.scala 115:36 connections.scala 50:12]
  wire [12:0] _GEN_88 = _T_54 ? {{7'd0}, _T_52} : _T_41; // @[Conditional.scala 39:67 Decode.scala 117:18 Decode.scala 72:12]
  wire  _GEN_89 = _T_54 | _T_44; // @[Conditional.scala 39:67 Decode.scala 118:22]
  wire  _GEN_90 = _T_53 & dual; // @[Conditional.scala 39:67 Decode.scala 110:36 connections.scala 49:12]
  wire  _GEN_91 = _T_53 | _GEN_89; // @[Conditional.scala 39:67 Decode.scala 111:22]
  wire  _GEN_92 = _T_53 ? _GEN_82 : _GEN_85; // @[Conditional.scala 39:67]
  wire  _GEN_93 = _T_53 ? 1'h0 : _GEN_86; // @[Conditional.scala 39:67 connections.scala 50:12]
  wire [12:0] _GEN_95 = _T_53 ? _T_41 : _GEN_88; // @[Conditional.scala 39:67 Decode.scala 72:12]
  wire  _GEN_96 = _T_51 & dual; // @[Conditional.scala 39:67 Decode.scala 104:35 connections.scala 48:11]
  wire  _GEN_97 = _T_51 ? dual : _GEN_92; // @[Conditional.scala 39:67 Decode.scala 105:29]
  wire [12:0] _GEN_98 = _T_51 ? {{7'd0}, _T_52} : _GEN_95; // @[Conditional.scala 39:67 Decode.scala 106:18]
  wire  _GEN_99 = _T_51 | _GEN_91; // @[Conditional.scala 39:67 Decode.scala 107:22]
  wire  _GEN_100 = _T_51 ? 1'h0 : _GEN_90; // @[Conditional.scala 39:67 connections.scala 49:12]
  wire  _GEN_101 = _T_51 ? _GEN_82 : _GEN_92; // @[Conditional.scala 39:67]
  wire  _GEN_102 = _T_51 ? 1'h0 : _GEN_93; // @[Conditional.scala 39:67 connections.scala 50:12]
  wire  _GEN_103 = _T_50 ? dual : _GEN_96; // @[Conditional.scala 39:67 Decode.scala 100:35]
  wire  _GEN_104 = _T_50 | _GEN_99; // @[Conditional.scala 39:67 Decode.scala 101:22]
  wire  _GEN_105 = _T_50 ? _GEN_82 : _GEN_97; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_106 = _T_50 ? _T_41 : _GEN_98; // @[Conditional.scala 39:67 Decode.scala 72:12]
  wire  _GEN_107 = _T_50 ? 1'h0 : _GEN_100; // @[Conditional.scala 39:67 connections.scala 49:12]
  wire  _GEN_108 = _T_50 ? _GEN_82 : _GEN_101; // @[Conditional.scala 39:67]
  wire  _GEN_109 = _T_50 ? 1'h0 : _GEN_102; // @[Conditional.scala 39:67 connections.scala 50:12]
  wire  _GEN_110 = _T_49 & dual; // @[Conditional.scala 39:67 Decode.scala 96:35 connections.scala 47:11]
  wire  _GEN_111 = _T_49 | _GEN_104; // @[Conditional.scala 39:67 Decode.scala 97:22]
  wire  _GEN_112 = _T_49 ? 1'h0 : _GEN_103; // @[Conditional.scala 39:67 connections.scala 48:11]
  wire  _GEN_113 = _T_49 ? _GEN_82 : _GEN_105; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_114 = _T_49 ? _T_41 : _GEN_106; // @[Conditional.scala 39:67 Decode.scala 72:12]
  wire  _GEN_115 = _T_49 ? 1'h0 : _GEN_107; // @[Conditional.scala 39:67 connections.scala 49:12]
  wire  _GEN_116 = _T_49 ? _GEN_82 : _GEN_108; // @[Conditional.scala 39:67]
  wire  _GEN_117 = _T_49 ? 1'h0 : _GEN_109; // @[Conditional.scala 39:67 connections.scala 50:12]
  wire  _GEN_118 = _T_48 ? dual : _GEN_116; // @[Conditional.scala 39:67 Decode.scala 92:28]
  wire  _GEN_119 = _T_48 | _GEN_111; // @[Conditional.scala 39:67 Decode.scala 93:22]
  wire  _GEN_121 = _T_48 ? 1'h0 : _GEN_112; // @[Conditional.scala 39:67 connections.scala 48:11]
  wire  _GEN_122 = _T_48 ? _GEN_82 : _GEN_113; // @[Conditional.scala 39:67]
  wire [12:0] _GEN_123 = _T_48 ? _T_41 : _GEN_114; // @[Conditional.scala 39:67 Decode.scala 72:12]
  wire  _GEN_124 = _T_48 ? 1'h0 : _GEN_115; // @[Conditional.scala 39:67 connections.scala 49:12]
  wire  _GEN_125 = _T_48 ? 1'h0 : _GEN_117; // @[Conditional.scala 39:67 connections.scala 50:12]
  wire  _GEN_126 = _T_47 ? dual : _GEN_118; // @[Conditional.scala 40:58 Decode.scala 88:28]
  wire  _GEN_127 = _T_47 | _GEN_119; // @[Conditional.scala 40:58 Decode.scala 89:22]
  wire  _GEN_129 = _T_47 ? 1'h0 : _GEN_121; // @[Conditional.scala 40:58 connections.scala 48:11]
  wire  _GEN_130 = _T_47 ? _GEN_82 : _GEN_122; // @[Conditional.scala 40:58]
  wire [12:0] _GEN_131 = _T_47 ? _T_41 : _GEN_123; // @[Conditional.scala 40:58 Decode.scala 72:12]
  wire  _GEN_132 = _T_47 ? 1'h0 : _GEN_124; // @[Conditional.scala 40:58 connections.scala 49:12]
  wire  _GEN_133 = _T_47 ? 1'h0 : _GEN_125; // @[Conditional.scala 40:58 connections.scala 50:12]
  wire  _GEN_134 = decReg_instr_b[26:22] == 5'h8 ? _GEN_126 : _GEN_82; // @[Decode.scala 85:33]
  wire  _GEN_135 = decReg_instr_b[26:22] == 5'h8 ? _GEN_127 : _T_44; // @[Decode.scala 85:33]
  wire  _GEN_137 = decReg_instr_b[26:22] == 5'h8 & _GEN_129; // @[Decode.scala 85:33 connections.scala 48:11]
  wire  _GEN_138 = decReg_instr_b[26:22] == 5'h8 ? _GEN_130 : _GEN_82; // @[Decode.scala 85:33]
  wire [12:0] _GEN_139 = decReg_instr_b[26:22] == 5'h8 ? _GEN_131 : _T_41; // @[Decode.scala 85:33 Decode.scala 72:12]
  wire  _GEN_140 = decReg_instr_b[26:22] == 5'h8 & _GEN_132; // @[Decode.scala 85:33 connections.scala 49:12]
  wire  _GEN_141 = decReg_instr_b[26:22] == 5'h8 & _GEN_133; // @[Decode.scala 85:33 connections.scala 50:12]
  wire  _GEN_142 = _T_50 & dual; // @[Conditional.scala 39:67 Decode.scala 130:35 connections.scala 52:11]
  wire  _GEN_143 = _T_50 ? dual : _GEN_134; // @[Conditional.scala 39:67 Decode.scala 131:28]
  wire  _GEN_144 = _T_50 | _GEN_135; // @[Conditional.scala 39:67 Decode.scala 132:22]
  wire  _GEN_146 = _T_49 | _GEN_144; // @[Conditional.scala 40:58 Decode.scala 127:22]
  wire  _GEN_147 = _T_49 ? 1'h0 : _GEN_142; // @[Conditional.scala 40:58 connections.scala 52:11]
  wire  _GEN_148 = _T_49 ? _GEN_134 : _GEN_143; // @[Conditional.scala 40:58]
  wire  _GEN_149 = decReg_instr_b[26:22] == 5'h9 & _GEN_110; // @[Decode.scala 123:33 connections.scala 51:11]
  wire  decoded_1 = decReg_instr_b[26:22] == 5'h9 ? _GEN_146 : _GEN_135; // @[Decode.scala 123:33]
  wire  _GEN_151 = decReg_instr_b[26:22] == 5'h9 & _GEN_147; // @[Decode.scala 123:33 connections.scala 52:11]
  wire  _GEN_152 = decReg_instr_b[26:22] == 5'h9 ? _GEN_148 : _GEN_134; // @[Decode.scala 123:33]
  wire  hi_1 = decReg_instr_b[3]; // @[Decode.scala 141:41]
  wire  lo_9 = decReg_instr_b[0]; // @[Decode.scala 141:51]
  wire [1:0] _T_59 = {hi_1,lo_9}; // @[Cat.scala 30:58]
  wire [2:0] ldsize = decReg_instr_a[11:9]; // @[Decode.scala 156:21]
  wire [1:0] ldtype = decReg_instr_a[8:7]; // @[Decode.scala 157:21]
  wire [2:0] stsize = decReg_instr_a[21:19]; // @[Decode.scala 158:21]
  wire [1:0] sttype = decReg_instr_a[18:17]; // @[Decode.scala 159:21]
  wire [3:0] stcfun = decReg_instr_a[21:18]; // @[Decode.scala 160:21]
  wire [17:0] hi_lo = decReg_instr_a[17:0]; // @[Decode.scala 169:34]
  wire [20:0] stcImm = {1'h0,hi_lo,2'h0}; // @[Cat.scala 30:58]
  wire  longImm = decReg_instr_a[26:22] == 5'h1f & decReg_instr_a[6:4] == 3'h0; // @[Decode.scala 183:31]
  wire [3:0] _GEN_153 = longImm ? decReg_instr_a[3:0] : _GEN_9; // @[Decode.scala 183:59 Decode.scala 184:28]
  wire  _GEN_154 = longImm | _GEN_66; // @[Decode.scala 183:59 Decode.scala 185:23]
  wire  _GEN_156 = longImm | _GEN_80; // @[Decode.scala 183:59 Decode.scala 187:22]
  wire  _GEN_157 = longImm | _GEN_78; // @[Decode.scala 183:59 Decode.scala 188:16]
  wire  _T_71 = 4'h0 == stcfun; // @[Conditional.scala 37:30]
  wire  _T_72 = 4'h4 == stcfun; // @[Conditional.scala 37:30]
  wire  _T_73 = 4'h5 == stcfun; // @[Conditional.scala 37:30]
  wire  _T_74 = 4'h8 == stcfun; // @[Conditional.scala 37:30]
  wire  _T_75 = 4'hc == stcfun; // @[Conditional.scala 37:30]
  wire  _T_76 = 4'hd == stcfun; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_159 = _T_76 ? 3'h6 : 3'h0; // @[Conditional.scala 39:67 Decode.scala 224:26 connections.scala 146:13]
  wire  _GEN_160 = _T_76 | _GEN_157; // @[Conditional.scala 39:67 Decode.scala 225:20]
  wire  _GEN_161 = _T_75 | _T_76; // @[Conditional.scala 39:67 Decode.scala 217:15]
  wire [2:0] _GEN_162 = _T_75 ? 3'h6 : _GEN_159; // @[Conditional.scala 39:67 Decode.scala 218:26]
  wire  _GEN_163 = _T_75 | _GEN_154; // @[Conditional.scala 39:67 Decode.scala 219:27]
  wire  _GEN_164 = _T_75 | _GEN_160; // @[Conditional.scala 39:67 Decode.scala 220:20]
  wire  _GEN_165 = _T_74 | _GEN_161; // @[Conditional.scala 39:67 Decode.scala 211:15]
  wire [2:0] _GEN_166 = _T_74 ? 3'h5 : _GEN_162; // @[Conditional.scala 39:67 Decode.scala 212:26]
  wire  _GEN_167 = _T_74 | _GEN_163; // @[Conditional.scala 39:67 Decode.scala 213:27]
  wire  _GEN_168 = _T_74 | _GEN_164; // @[Conditional.scala 39:67 Decode.scala 214:20]
  wire  _GEN_169 = _T_73 | _GEN_165; // @[Conditional.scala 39:67 Decode.scala 206:15]
  wire [2:0] _GEN_170 = _T_73 ? 3'h4 : _GEN_166; // @[Conditional.scala 39:67 Decode.scala 207:26]
  wire  _GEN_171 = _T_73 | _GEN_168; // @[Conditional.scala 39:67 Decode.scala 208:20]
  wire  _GEN_172 = _T_73 ? _GEN_154 : _GEN_167; // @[Conditional.scala 39:67]
  wire  _GEN_173 = _T_72 | _GEN_169; // @[Conditional.scala 39:67 Decode.scala 200:15]
  wire [2:0] _GEN_174 = _T_72 ? 3'h4 : _GEN_170; // @[Conditional.scala 39:67 Decode.scala 201:26]
  wire  _GEN_175 = _T_72 | _GEN_172; // @[Conditional.scala 39:67 Decode.scala 202:27]
  wire  _GEN_176 = _T_72 | _GEN_171; // @[Conditional.scala 39:67 Decode.scala 203:20]
  wire  _GEN_177 = _T_71 | _GEN_173; // @[Conditional.scala 40:58 Decode.scala 194:15]
  wire [2:0] _GEN_178 = _T_71 ? 3'h3 : _GEN_174; // @[Conditional.scala 40:58 Decode.scala 195:26]
  wire  _GEN_179 = _T_71 | _GEN_175; // @[Conditional.scala 40:58 Decode.scala 196:27]
  wire  _GEN_180 = _T_71 | _GEN_176; // @[Conditional.scala 40:58 Decode.scala 197:20]
  wire  isSTC = decReg_instr_a[26:22] == 5'hc & _GEN_177; // @[Decode.scala 191:31 Decode.scala 177:9]
  wire [2:0] _GEN_182 = decReg_instr_a[26:22] == 5'hc ? _GEN_178 : 3'h0; // @[Decode.scala 191:31 connections.scala 146:13]
  wire  _GEN_183 = decReg_instr_a[26:22] == 5'hc ? _GEN_179 : _GEN_154; // @[Decode.scala 191:31]
  wire  _GEN_184 = decReg_instr_a[26:22] == 5'hc ? _GEN_180 : _GEN_157; // @[Decode.scala 191:31]
  wire  _T_77 = decReg_instr_a[26:22] == 5'h16; // @[Decode.scala 231:15]
  wire [4:0] _GEN_186 = decReg_instr_a[26:22] == 5'h16 ? decReg_instr_a[4:0] : 5'h0; // @[Decode.scala 231:36 Decode.scala 233:19 connections.scala 160:10]
  wire  _GEN_187 = decReg_instr_a[26:22] == 5'h16 | _GEN_184; // @[Decode.scala 231:36 Decode.scala 234:16]
  wire  _T_81 = decReg_instr_a[26:22] == 5'h11 | decReg_instr_a[26:22] == 5'h10; // @[Decode.scala 236:35]
  wire  _GEN_188 = decReg_instr_a[26:22] == 5'h11 | decReg_instr_a[26:22] == 5'h10 | _GEN_183; // @[Decode.scala 236:68 Decode.scala 237:23]
  wire  _GEN_190 = (decReg_instr_a[26:22] == 5'h11 | decReg_instr_a[26:22] == 5'h10) & decReg_instr_a[26:22] == 5'h10; // @[Decode.scala 236:68 Decode.scala 239:25 connections.scala 161:16]
  wire  _GEN_191 = decReg_instr_a[26:22] == 5'h11 | decReg_instr_a[26:22] == 5'h10 | _GEN_187; // @[Decode.scala 236:68 Decode.scala 240:16]
  wire  _T_85 = decReg_instr_a[26:22] == 5'h13 | decReg_instr_a[26:22] == 5'h12; // @[Decode.scala 242:33]
  wire  _GEN_192 = decReg_instr_a[26:22] == 5'h13 | decReg_instr_a[26:22] == 5'h12 | _GEN_188; // @[Decode.scala 242:64 Decode.scala 243:23]
  wire  _GEN_194 = decReg_instr_a[26:22] == 5'h13 | decReg_instr_a[26:22] == 5'h12 ? decReg_instr_a[26:22] == 5'h12 :
    _GEN_190; // @[Decode.scala 242:64 Decode.scala 245:25]
  wire  _GEN_195 = decReg_instr_a[26:22] == 5'h13 | decReg_instr_a[26:22] == 5'h12 | _GEN_191; // @[Decode.scala 242:64 Decode.scala 246:16]
  wire  _T_89 = decReg_instr_a[26:22] == 5'h15 | decReg_instr_a[26:22] == 5'h14; // @[Decode.scala 248:35]
  wire  _GEN_196 = decReg_instr_a[26:22] == 5'h15 | decReg_instr_a[26:22] == 5'h14 | _GEN_192; // @[Decode.scala 248:68 Decode.scala 249:23]
  wire  _GEN_198 = decReg_instr_a[26:22] == 5'h15 | decReg_instr_a[26:22] == 5'h14 ? decReg_instr_a[26:22] == 5'h14 :
    _GEN_194; // @[Decode.scala 248:68 Decode.scala 251:25]
  wire  _GEN_199 = decReg_instr_a[26:22] == 5'h15 | decReg_instr_a[26:22] == 5'h14 | _GEN_195; // @[Decode.scala 248:68 Decode.scala 252:16]
  wire  _T_94 = 4'h0 == decReg_instr_a[3:0]; // @[Conditional.scala 37:30]
  wire  _T_95 = 4'h1 == decReg_instr_a[3:0]; // @[Conditional.scala 37:30]
  wire  _T_96 = 4'h4 == decReg_instr_a[3:0]; // @[Conditional.scala 37:30]
  wire  _T_97 = 4'h5 == decReg_instr_a[3:0]; // @[Conditional.scala 37:30]
  wire  _T_98 = 4'ha == decReg_instr_a[3:0]; // @[Conditional.scala 37:30]
  wire  _GEN_200 = _T_98 | _T_89; // @[Conditional.scala 39:67 Decode.scala 273:23]
  wire  _GEN_201 = _T_98 | _GEN_199; // @[Conditional.scala 39:67 Decode.scala 274:20]
  wire  _GEN_202 = _T_97 | _T_85; // @[Conditional.scala 39:67 Decode.scala 269:31]
  wire  _GEN_203 = _T_97 | _GEN_201; // @[Conditional.scala 39:67 Decode.scala 270:20]
  wire  _GEN_204 = _T_97 ? _T_89 : _GEN_200; // @[Conditional.scala 39:67]
  wire  _GEN_205 = _T_96 | _T_81; // @[Conditional.scala 39:67 Decode.scala 265:23]
  wire  _GEN_206 = _T_96 | _GEN_203; // @[Conditional.scala 39:67 Decode.scala 266:20]
  wire  _GEN_207 = _T_96 ? _T_85 : _GEN_202; // @[Conditional.scala 39:67]
  wire  _GEN_208 = _T_96 ? _T_89 : _GEN_204; // @[Conditional.scala 39:67]
  wire  _GEN_210 = _T_95 | _GEN_206; // @[Conditional.scala 39:67 Decode.scala 262:20]
  wire  _GEN_211 = _T_95 ? _T_81 : _GEN_205; // @[Conditional.scala 39:67]
  wire  _GEN_212 = _T_95 ? _T_85 : _GEN_207; // @[Conditional.scala 39:67]
  wire  _GEN_213 = _T_95 ? _T_89 : _GEN_208; // @[Conditional.scala 39:67]
  wire  _GEN_215 = _T_94 | _GEN_210; // @[Conditional.scala 40:58 Decode.scala 258:20]
  wire  _GEN_216 = _T_94 ? 1'h0 : _T_95; // @[Conditional.scala 40:58 connections.scala 159:10]
  wire  _GEN_217 = _T_94 ? _T_81 : _GEN_211; // @[Conditional.scala 40:58]
  wire  _GEN_218 = _T_94 ? _T_85 : _GEN_212; // @[Conditional.scala 40:58]
  wire  _GEN_219 = _T_94 ? _T_89 : _GEN_213; // @[Conditional.scala 40:58]
  wire  _GEN_220 = (decReg_instr_a[26:22] == 5'h19 | decReg_instr_a[26:22] == 5'h18) & _T_94; // @[Decode.scala 254:68 connections.scala 155:9]
  wire  _GEN_221 = decReg_instr_a[26:22] == 5'h19 | decReg_instr_a[26:22] == 5'h18 ? _GEN_215 : _GEN_199; // @[Decode.scala 254:68]
  wire  _GEN_222 = (decReg_instr_a[26:22] == 5'h19 | decReg_instr_a[26:22] == 5'h18) & _GEN_216; // @[Decode.scala 254:68 connections.scala 159:10]
  wire  _GEN_223 = decReg_instr_a[26:22] == 5'h19 | decReg_instr_a[26:22] == 5'h18 ? _GEN_217 : _T_81; // @[Decode.scala 254:68]
  wire  _GEN_224 = decReg_instr_a[26:22] == 5'h19 | decReg_instr_a[26:22] == 5'h18 ? _GEN_218 : _T_85; // @[Decode.scala 254:68]
  wire  _GEN_225 = decReg_instr_a[26:22] == 5'h19 | decReg_instr_a[26:22] == 5'h18 ? _GEN_219 : _T_89; // @[Decode.scala 254:68]
  wire  _GEN_226 = decReg_instr_a[26:22] == 5'h19 | decReg_instr_a[26:22] == 5'h18 ? decReg_instr_a[26:22] == 5'h18 :
    _GEN_198; // @[Decode.scala 254:68 Decode.scala 277:25]
  wire  _T_100 = decReg_instr_a[26:22] == 5'ha; // @[Decode.scala 283:15]
  wire  _T_101 = 3'h0 == ldsize; // @[Conditional.scala 37:30]
  wire  _T_102 = 3'h1 == ldsize; // @[Conditional.scala 37:30]
  wire  _T_103 = 3'h2 == ldsize; // @[Conditional.scala 37:30]
  wire  _T_104 = 3'h3 == ldsize; // @[Conditional.scala 37:30]
  wire  _T_105 = 3'h4 == ldsize; // @[Conditional.scala 37:30]
  wire  _GEN_229 = _T_104 | _T_105; // @[Conditional.scala 39:67 Decode.scala 301:29]
  wire  _GEN_230 = _T_104 ? 1'h0 : _T_105; // @[Conditional.scala 39:67 connections.scala 94:10]
  wire  _GEN_231 = _T_103 | _GEN_230; // @[Conditional.scala 39:67 Decode.scala 296:29]
  wire  _GEN_232 = _T_103 ? 1'h0 : _T_104; // @[Conditional.scala 39:67 Decode.scala 281:9]
  wire  _GEN_233 = _T_103 ? 1'h0 : _GEN_229; // @[Conditional.scala 39:67 connections.scala 95:10]
  wire  _GEN_234 = _T_102 | _GEN_232; // @[Conditional.scala 39:67 Decode.scala 292:15]
  wire  _GEN_235 = _T_102 ? 1'h0 : _GEN_231; // @[Conditional.scala 39:67 connections.scala 94:10]
  wire  _GEN_236 = _T_102 ? 1'h0 : _GEN_233; // @[Conditional.scala 39:67 connections.scala 95:10]
  wire [1:0] _GEN_237 = _T_101 ? 2'h2 : {{1'd0}, _GEN_234}; // @[Conditional.scala 40:58 Decode.scala 289:15]
  wire  _GEN_238 = _T_101 ? 1'h0 : _GEN_234; // @[Conditional.scala 40:58 connections.scala 93:11]
  wire  _GEN_239 = _T_101 ? 1'h0 : _GEN_235; // @[Conditional.scala 40:58 connections.scala 94:10]
  wire  _GEN_240 = _T_101 ? 1'h0 : _GEN_236; // @[Conditional.scala 40:58 connections.scala 95:10]
  wire [1:0] _GEN_241 = ldtype == 2'h2 & io_exc_local ? 2'h1 : ldtype; // @[Decode.scala 309:46 Decode.scala 310:26 Decode.scala 308:24]
  wire  _T_108 = ldtype == 2'h0; // @[Decode.scala 312:17]
  wire  _GEN_244 = decReg_instr_a[26:22] == 5'ha | _GEN_156; // @[Decode.scala 283:31 Decode.scala 286:22]
  wire [1:0] _GEN_245 = decReg_instr_a[26:22] == 5'ha ? _GEN_237 : 2'h0; // @[Decode.scala 283:31 Decode.scala 281:9]
  wire  _GEN_246 = decReg_instr_a[26:22] == 5'ha & _GEN_238; // @[Decode.scala 283:31 connections.scala 93:11]
  wire  _GEN_247 = decReg_instr_a[26:22] == 5'ha & _GEN_239; // @[Decode.scala 283:31 connections.scala 94:10]
  wire  _GEN_248 = decReg_instr_a[26:22] == 5'ha & _GEN_240; // @[Decode.scala 283:31 connections.scala 95:10]
  wire [1:0] _GEN_249 = decReg_instr_a[26:22] == 5'ha ? _GEN_241 : 2'h0; // @[Decode.scala 283:31 connections.scala 96:9]
  wire  _GEN_250 = decReg_instr_a[26:22] == 5'ha & _T_108; // @[Decode.scala 283:31 Decode.scala 176:11]
  wire  _GEN_251 = decReg_instr_a[26:22] == 5'ha | _GEN_221; // @[Decode.scala 283:31 Decode.scala 315:16]
  wire  _T_109 = decReg_instr_a[26:22] == 5'hb; // @[Decode.scala 318:15]
  wire  _T_110 = 3'h0 == stsize; // @[Conditional.scala 37:30]
  wire  _T_111 = 3'h1 == stsize; // @[Conditional.scala 37:30]
  wire  _T_112 = 3'h2 == stsize; // @[Conditional.scala 37:30]
  wire  _GEN_252 = _T_112 | _GEN_247; // @[Conditional.scala 39:67 Decode.scala 330:29]
  wire [1:0] _GEN_253 = _T_111 ? 2'h1 : _GEN_245; // @[Conditional.scala 39:67 Decode.scala 326:15]
  wire  _GEN_254 = _T_111 | _GEN_246; // @[Conditional.scala 39:67 Decode.scala 327:30]
  wire  _GEN_255 = _T_111 ? _GEN_247 : _GEN_252; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_256 = _T_110 ? 2'h2 : _GEN_253; // @[Conditional.scala 40:58 Decode.scala 323:15]
  wire  _GEN_257 = _T_110 ? _GEN_246 : _GEN_254; // @[Conditional.scala 40:58]
  wire  _GEN_258 = _T_110 ? _GEN_247 : _GEN_255; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_259 = sttype == 2'h2 & io_exc_local ? 2'h1 : sttype; // @[Decode.scala 334:46 Decode.scala 335:26 Decode.scala 333:24]
  wire  _GEN_260 = sttype == 2'h0 | _GEN_250; // @[Decode.scala 337:30 Decode.scala 338:15]
  wire  isMem = decReg_instr_a[26:22] == 5'hb | _T_100; // @[Decode.scala 318:31 Decode.scala 319:11]
  wire [1:0] shamt = decReg_instr_a[26:22] == 5'hb ? _GEN_256 : _GEN_245; // @[Decode.scala 318:31]
  wire  _GEN_264 = decReg_instr_a[26:22] == 5'hb ? _GEN_257 : _GEN_246; // @[Decode.scala 318:31]
  wire  _GEN_265 = decReg_instr_a[26:22] == 5'hb ? _GEN_258 : _GEN_247; // @[Decode.scala 318:31]
  wire [1:0] _GEN_266 = decReg_instr_a[26:22] == 5'hb ? _GEN_259 : _GEN_249; // @[Decode.scala 318:31]
  wire  isStack = decReg_instr_a[26:22] == 5'hb ? _GEN_260 : _GEN_250; // @[Decode.scala 318:31]
  wire  decoded_0 = decReg_instr_a[26:22] == 5'hb | _GEN_251; // @[Decode.scala 318:31 Decode.scala 340:16]
  wire [6:0] lo_10 = decReg_instr_a[6:0]; // @[Decode.scala 345:32]
  wire [7:0] _T_116 = {1'h0,lo_10}; // @[Cat.scala 30:58]
  wire  _T_117 = 2'h1 == shamt; // @[Conditional.scala 37:30]
  wire [8:0] _T_118 = {1'h0,lo_10,1'h0}; // @[Cat.scala 30:58]
  wire  _T_119 = 2'h2 == shamt; // @[Conditional.scala 37:30]
  wire [9:0] _T_120 = {1'h0,lo_10,2'h0}; // @[Cat.scala 30:58]
  wire [9:0] _GEN_269 = _T_119 ? _T_120 : {{2'd0}, _T_116}; // @[Conditional.scala 39:67 Decode.scala 348:27 Decode.scala 345:11]
  wire [9:0] addrImm = _T_117 ? {{1'd0}, _T_118} : _GEN_269; // @[Conditional.scala 40:58 Decode.scala 347:27]
  wire [31:0] _T_124 = isMem ? {{22'd0}, addrImm} : decReg_instr_b; // @[Decode.scala 355:38]
  wire [31:0] _T_125 = isStack ? {{22'd0}, addrImm} : _T_124; // @[Decode.scala 354:34]
  wire [31:0] _T_126 = isSTC ? {{11'd0}, stcImm} : _T_125; // @[Decode.scala 353:30]
  wire [31:0] _GEN_271 = isSTC | isStack | isMem | longImm ? _T_126 : {{19'd0}, _GEN_67}; // @[Decode.scala 352:47 Decode.scala 353:24 Decode.scala 138:24]
  wire [21:0] hi_lo_3 = decReg_instr_a[21:0]; // @[Decode.scala 361:42]
  wire [24:0] _T_127 = {1'h0,hi_lo_3,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] hi_6 = decReg_instr_a[21] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [29:0] _T_130 = {hi_6,hi_lo_3}; // @[Cat.scala 30:58]
  wire [29:0] _T_132 = decReg_pc + _T_130; // @[Decode.scala 365:38]
  wire  _GEN_272 = io_decex_rdAddr_0 == 5'h0 ? 1'h0 : _GEN_244; // @[Decode.scala 378:49 Decode.scala 379:24]
  wire  _GEN_273 = io_decex_rdAddr_1 == 5'h0 ? 1'h0 : _GEN_152; // @[Decode.scala 378:49 Decode.scala 379:24]
  wire  _T_136 = dual ? decoded_0 & decoded_1 : decoded_0; // @[Decode.scala 384:25]
  reg [1:0] inDelaySlot; // @[Decode.scala 387:24]
  wire  _T_139 = io_exc_intr & inDelaySlot == 2'h0; // @[Decode.scala 390:21]
  wire  _T_140 = io_exc_exc | _T_139; // @[Decode.scala 389:19]
  wire [29:0] _T_143 = io_exc_exc ? io_exc_excBase : decReg_base; // @[Decode.scala 397:25]
  wire [29:0] _T_144 = io_exc_exc ? io_exc_excAddr : decReg_relPc; // @[Decode.scala 398:26]
  wire [12:0] _GEN_321 = _T_140 ? 13'h0 : _GEN_139; // @[Decode.scala 390:50 connections.scala 150:12 Decode.scala 138:24]
  wire [1:0] _T_146 = inDelaySlot - 2'h1; // @[Decode.scala 403:36]
  wire  _T_149 = io_decex_call | io_decex_ret | io_decex_brcf | io_decex_xcall; // @[Decode.scala 405:75]
  wire  _T_150 = _T_149 | io_decex_xret; // @[Decode.scala 406:43]
  wire [1:0] _T_152 = inDelaySlot > 2'h1 ? _T_146 : 2'h1; // @[Decode.scala 409:39]
  wire [1:0] _T_154 = inDelaySlot != 2'h0 ? _T_146 : 2'h0; // @[Decode.scala 410:39]
  wire [1:0] _T_155 = io_decex_aluOp_0_isMul ? _T_152 : _T_154; // @[Decode.scala 408:35]
  RegisterFile rf ( // @[Decode.scala 19:18]
    .clock(rf_clock),
    .io_ena(rf_io_ena),
    .io_rfRead_rsAddr_0(rf_io_rfRead_rsAddr_0),
    .io_rfRead_rsAddr_1(rf_io_rfRead_rsAddr_1),
    .io_rfRead_rsAddr_2(rf_io_rfRead_rsAddr_2),
    .io_rfRead_rsAddr_3(rf_io_rfRead_rsAddr_3),
    .io_rfRead_rsData_0(rf_io_rfRead_rsData_0),
    .io_rfRead_rsData_1(rf_io_rfRead_rsData_1),
    .io_rfRead_rsData_2(rf_io_rfRead_rsData_2),
    .io_rfRead_rsData_3(rf_io_rfRead_rsData_3),
    .io_rfWrite_0_addr(rf_io_rfWrite_0_addr),
    .io_rfWrite_0_data(rf_io_rfWrite_0_data),
    .io_rfWrite_0_valid(rf_io_rfWrite_0_valid),
    .io_rfWrite_1_addr(rf_io_rfWrite_1_addr),
    .io_rfWrite_1_data(rf_io_rfWrite_1_data),
    .io_rfWrite_1_valid(rf_io_rfWrite_1_valid)
  );
  assign io_decex_base = _T_140 ? _T_143 : decReg_base; // @[Decode.scala 390:50 Decode.scala 397:19 Decode.scala 370:17]
  assign io_decex_relPc = _T_140 ? _T_144 : decReg_relPc; // @[Decode.scala 390:50 Decode.scala 398:20 Decode.scala 371:18]
  assign io_decex_pred_0 = _T_140 ? 4'h0 : decReg_instr_a[30:27]; // @[Decode.scala 390:50 Decode.scala 392:22 Decode.scala 145:22]
  assign io_decex_pred_1 = _T_140 ? 4'h8 : decReg_instr_b[30:27]; // @[Decode.scala 390:50 connections.scala 141:10 Decode.scala 145:22]
  assign io_decex_aluOp_0_func = _T_140 ? 4'h0 : _GEN_153; // @[Decode.scala 390:50 connections.scala 46:10]
  assign io_decex_aluOp_0_isMul = _T_140 ? 1'h0 : _GEN_64; // @[Decode.scala 390:50 connections.scala 47:11]
  assign io_decex_aluOp_0_isCmp = _T_140 ? 1'h0 : _GEN_65; // @[Decode.scala 390:50 connections.scala 48:11]
  assign io_decex_aluOp_0_isPred = _T_140 ? 1'h0 : _GEN_68; // @[Decode.scala 390:50 connections.scala 49:12]
  assign io_decex_aluOp_0_isBCpy = _T_140 ? 1'h0 : _GEN_69; // @[Decode.scala 390:50 connections.scala 50:12]
  assign io_decex_aluOp_0_isMTS = _T_140 ? 1'h0 : _GEN_77; // @[Decode.scala 390:50 connections.scala 51:11]
  assign io_decex_aluOp_0_isMFS = _T_140 ? 1'h0 : _GEN_79; // @[Decode.scala 390:50 connections.scala 52:11]
  assign io_decex_aluOp_1_func = _T_140 ? 4'h0 : _GEN_81; // @[Decode.scala 390:50 connections.scala 46:10]
  assign io_decex_aluOp_1_isCmp = _T_140 ? 1'h0 : _GEN_137; // @[Decode.scala 390:50 connections.scala 48:11]
  assign io_decex_aluOp_1_isPred = _T_140 ? 1'h0 : _GEN_140; // @[Decode.scala 390:50 connections.scala 49:12]
  assign io_decex_aluOp_1_isBCpy = _T_140 ? 1'h0 : _GEN_141; // @[Decode.scala 390:50 connections.scala 50:12]
  assign io_decex_aluOp_1_isMTS = _T_140 ? 1'h0 : _GEN_149; // @[Decode.scala 390:50 connections.scala 51:11]
  assign io_decex_aluOp_1_isMFS = _T_140 ? 1'h0 : _GEN_151; // @[Decode.scala 390:50 connections.scala 52:11]
  assign io_decex_predOp_0_func = _T_140 ? 2'h0 : _T_33; // @[Decode.scala 390:50 connections.scala 63:10 Decode.scala 141:29]
  assign io_decex_predOp_0_dest = _T_140 ? 3'h0 : decReg_instr_a[19:17]; // @[Decode.scala 390:50 connections.scala 64:10 Decode.scala 144:29]
  assign io_decex_predOp_0_s1Addr = _T_140 ? 4'h0 : decReg_instr_a[15:12]; // @[Decode.scala 390:50 connections.scala 65:12 Decode.scala 142:31]
  assign io_decex_predOp_0_s2Addr = _T_140 ? 4'h0 : decReg_instr_a[10:7]; // @[Decode.scala 390:50 connections.scala 66:12 Decode.scala 143:31]
  assign io_decex_predOp_1_func = _T_140 ? 2'h0 : _T_59; // @[Decode.scala 390:50 connections.scala 63:10 Decode.scala 141:29]
  assign io_decex_predOp_1_dest = _T_140 ? 3'h0 : decReg_instr_b[19:17]; // @[Decode.scala 390:50 connections.scala 64:10 Decode.scala 144:29]
  assign io_decex_predOp_1_s1Addr = _T_140 ? 4'h0 : decReg_instr_b[15:12]; // @[Decode.scala 390:50 connections.scala 65:12 Decode.scala 142:31]
  assign io_decex_predOp_1_s2Addr = _T_140 ? 4'h0 : decReg_instr_b[10:7]; // @[Decode.scala 390:50 connections.scala 66:12 Decode.scala 143:31]
  assign io_decex_jmpOp_branch = _T_140 ? 1'h0 : _GEN_224; // @[Decode.scala 390:50 connections.scala 76:12]
  assign io_decex_jmpOp_target = _T_140 ? 30'h0 : _T_132; // @[Decode.scala 390:50 connections.scala 77:12 Decode.scala 365:25]
  assign io_decex_jmpOp_reloc = _T_140 ? 32'h0 : decReg_reloc; // @[Decode.scala 390:50 connections.scala 78:11 Decode.scala 366:24]
  assign io_decex_memOp_load = _T_140 ? 1'h0 : _T_100; // @[Decode.scala 390:50 connections.scala 91:10]
  assign io_decex_memOp_store = _T_140 ? 1'h0 : _T_109; // @[Decode.scala 390:50 connections.scala 92:11]
  assign io_decex_memOp_hword = _T_140 ? 1'h0 : _GEN_264; // @[Decode.scala 390:50 connections.scala 93:11]
  assign io_decex_memOp_byte = _T_140 ? 1'h0 : _GEN_265; // @[Decode.scala 390:50 connections.scala 94:10]
  assign io_decex_memOp_zext = _T_140 ? 1'h0 : _GEN_248; // @[Decode.scala 390:50 connections.scala 95:10]
  assign io_decex_memOp_typ = _T_140 ? 2'h0 : _GEN_266; // @[Decode.scala 390:50 connections.scala 96:9]
  assign io_decex_stackOp = _T_140 ? 3'h0 : _GEN_182; // @[Decode.scala 390:50 connections.scala 146:13]
  assign io_decex_rsAddr_0 = _T_140 ? 5'h0 : decReg_instr_a[16:12]; // @[Decode.scala 390:50 connections.scala 147:12 Decode.scala 45:22]
  assign io_decex_rsAddr_1 = _T_140 ? 5'h0 : decReg_instr_a[11:7]; // @[Decode.scala 390:50 connections.scala 147:12 Decode.scala 46:22]
  assign io_decex_rsAddr_2 = _T_140 ? 5'h0 : decReg_instr_b[16:12]; // @[Decode.scala 390:50 connections.scala 147:12 Decode.scala 48:24]
  assign io_decex_rsAddr_3 = _T_140 ? 5'h0 : decReg_instr_b[11:7]; // @[Decode.scala 390:50 connections.scala 147:12 Decode.scala 49:24]
  assign io_decex_rsData_0 = _T_140 ? 32'h0 : rf_io_rfRead_rsData_0; // @[Decode.scala 390:50 connections.scala 148:12 Decode.scala 52:22]
  assign io_decex_rsData_1 = _T_140 ? 32'h0 : rf_io_rfRead_rsData_1; // @[Decode.scala 390:50 connections.scala 148:12 Decode.scala 53:22]
  assign io_decex_rsData_2 = _T_140 ? 32'h0 : rf_io_rfRead_rsData_2; // @[Decode.scala 390:50 connections.scala 148:12 Decode.scala 55:24]
  assign io_decex_rsData_3 = _T_140 ? 32'h0 : rf_io_rfRead_rsData_3; // @[Decode.scala 390:50 connections.scala 148:12 Decode.scala 56:24]
  assign io_decex_rdAddr_0 = _T_140 ? 5'h0 : decReg_instr_a[21:17]; // @[Decode.scala 390:50 connections.scala 149:12 Decode.scala 374:22]
  assign io_decex_rdAddr_1 = _T_140 ? 5'h0 : decReg_instr_b[21:17]; // @[Decode.scala 390:50 connections.scala 149:12 Decode.scala 148:24]
  assign io_decex_immVal_0 = _T_140 ? 32'h0 : _GEN_271; // @[Decode.scala 390:50 connections.scala 150:12]
  assign io_decex_immVal_1 = {{19'd0}, _GEN_321}; // @[Decode.scala 390:50 connections.scala 150:12 Decode.scala 138:24]
  assign io_decex_immOp_0 = _T_140 | _GEN_196; // @[Decode.scala 390:50 Decode.scala 396:23]
  assign io_decex_immOp_1 = _T_140 ? 1'h0 : _GEN_138; // @[Decode.scala 390:50 connections.scala 151:11]
  assign io_decex_wrRd_0 = _T_140 ? 1'h0 : _GEN_272; // @[Decode.scala 390:50 connections.scala 152:10]
  assign io_decex_wrRd_1 = _T_140 ? 1'h0 : _GEN_273; // @[Decode.scala 390:50 connections.scala 152:10]
  assign io_decex_callAddr = _T_140 ? io_exc_addr : {{7'd0}, _T_127}; // @[Decode.scala 390:50 Decode.scala 395:23 Decode.scala 361:21]
  assign io_decex_call = _T_140 ? 1'h0 : _GEN_223; // @[Decode.scala 390:50 connections.scala 154:10]
  assign io_decex_ret = _T_140 ? 1'h0 : _GEN_220; // @[Decode.scala 390:50 connections.scala 155:9]
  assign io_decex_brcf = _T_140 ? 1'h0 : _GEN_225; // @[Decode.scala 390:50 connections.scala 156:10]
  assign io_decex_trap = _T_140 ? 1'h0 : _T_77; // @[Decode.scala 390:50 connections.scala 157:10]
  assign io_decex_xcall = io_exc_exc | _T_139; // @[Decode.scala 389:19]
  assign io_decex_xret = _T_140 ? 1'h0 : _GEN_222; // @[Decode.scala 390:50 connections.scala 159:10]
  assign io_decex_xsrc = _T_140 ? io_exc_src : _GEN_186; // @[Decode.scala 390:50 Decode.scala 394:19]
  assign io_decex_nonDelayed = _T_140 ? 1'h0 : _GEN_226; // @[Decode.scala 390:50 connections.scala 161:16]
  assign io_decex_illOp = _T_140 ? 1'h0 : ~_T_136; // @[Decode.scala 390:50 connections.scala 162:11 Decode.scala 384:18]
  assign rf_clock = clock;
  assign rf_io_ena = io_ena; // @[Decode.scala 27:13]
  assign rf_io_rfRead_rsAddr_0 = io_fedec_instr_a[16:12]; // @[Decode.scala 21:45]
  assign rf_io_rfRead_rsAddr_1 = io_fedec_instr_a[11:7]; // @[Decode.scala 22:45]
  assign rf_io_rfRead_rsAddr_2 = io_fedec_instr_b[16:12]; // @[Decode.scala 24:47]
  assign rf_io_rfRead_rsAddr_3 = io_fedec_instr_b[11:7]; // @[Decode.scala 25:47]
  assign rf_io_rfWrite_0_addr = io_rfWrite_0_addr; // @[Decode.scala 29:17]
  assign rf_io_rfWrite_0_data = io_rfWrite_0_data; // @[Decode.scala 29:17]
  assign rf_io_rfWrite_0_valid = io_rfWrite_0_valid; // @[Decode.scala 29:17]
  assign rf_io_rfWrite_1_addr = io_rfWrite_1_addr; // @[Decode.scala 29:17]
  assign rf_io_rfWrite_1_data = io_rfWrite_1_data; // @[Decode.scala 29:17]
  assign rf_io_rfWrite_1_valid = io_rfWrite_1_valid; // @[Decode.scala 29:17]
  always @(posedge clock) begin
    if (reset) begin // @[Decode.scala 414:15]
      decReg_instr_a <= 32'h0; // @[connections.scala 31:13]
    end else if (io_ena) begin // @[Decode.scala 33:16]
      if (io_flush) begin // @[Decode.scala 35:20]
        decReg_instr_a <= 32'h0; // @[connections.scala 31:13]
      end else begin
        decReg_instr_a <= io_fedec_instr_a; // @[Decode.scala 34:12]
      end
    end
    if (reset) begin // @[Decode.scala 414:15]
      decReg_instr_b <= 32'h0; // @[connections.scala 32:13]
    end else if (io_ena) begin // @[Decode.scala 33:16]
      if (io_flush) begin // @[Decode.scala 35:20]
        decReg_instr_b <= 32'h0; // @[connections.scala 32:13]
      end else begin
        decReg_instr_b <= io_fedec_instr_b; // @[Decode.scala 34:12]
      end
    end
    if (io_ena) begin // @[Decode.scala 33:16]
      decReg_pc <= io_fedec_pc; // @[Decode.scala 34:12]
    end
    if (io_ena) begin // @[Decode.scala 33:16]
      decReg_base <= io_fedec_base; // @[Decode.scala 34:12]
    end
    if (io_ena) begin // @[Decode.scala 33:16]
      decReg_reloc <= io_fedec_reloc; // @[Decode.scala 34:12]
    end
    if (io_ena) begin // @[Decode.scala 33:16]
      decReg_relPc <= io_fedec_relPc;
    end
    if (io_ena) begin // @[Decode.scala 402:16]
      if (io_flush) begin // @[Decode.scala 404:23]
        inDelaySlot <= 2'h1;
      end else if (_T_150) begin // @[Decode.scala 405:27]
        inDelaySlot <= 2'h3;
      end else if (io_decex_jmpOp_branch) begin // @[Decode.scala 407:31]
        inDelaySlot <= 2'h2;
      end else begin
        inDelaySlot <= _T_155;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  decReg_instr_a = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  decReg_instr_b = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  decReg_pc = _RAND_2[29:0];
  _RAND_3 = {1{`RANDOM}};
  decReg_base = _RAND_3[29:0];
  _RAND_4 = {1{`RANDOM}};
  decReg_reloc = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  decReg_relPc = _RAND_5[29:0];
  _RAND_6 = {1{`RANDOM}};
  inDelaySlot = _RAND_6[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Execute(
  input         clock,
  input         reset,
  input         io_ena,
  input         io_flush,
  output        io_brflush,
  input  [29:0] io_decex_base,
  input  [29:0] io_decex_relPc,
  input  [3:0]  io_decex_pred_0,
  input  [3:0]  io_decex_pred_1,
  input  [3:0]  io_decex_aluOp_0_func,
  input         io_decex_aluOp_0_isMul,
  input         io_decex_aluOp_0_isCmp,
  input         io_decex_aluOp_0_isPred,
  input         io_decex_aluOp_0_isBCpy,
  input         io_decex_aluOp_0_isMTS,
  input         io_decex_aluOp_0_isMFS,
  input  [3:0]  io_decex_aluOp_1_func,
  input         io_decex_aluOp_1_isCmp,
  input         io_decex_aluOp_1_isPred,
  input         io_decex_aluOp_1_isBCpy,
  input         io_decex_aluOp_1_isMTS,
  input         io_decex_aluOp_1_isMFS,
  input  [1:0]  io_decex_predOp_0_func,
  input  [2:0]  io_decex_predOp_0_dest,
  input  [3:0]  io_decex_predOp_0_s1Addr,
  input  [3:0]  io_decex_predOp_0_s2Addr,
  input  [1:0]  io_decex_predOp_1_func,
  input  [2:0]  io_decex_predOp_1_dest,
  input  [3:0]  io_decex_predOp_1_s1Addr,
  input  [3:0]  io_decex_predOp_1_s2Addr,
  input         io_decex_jmpOp_branch,
  input  [29:0] io_decex_jmpOp_target,
  input  [31:0] io_decex_jmpOp_reloc,
  input         io_decex_memOp_load,
  input         io_decex_memOp_store,
  input         io_decex_memOp_hword,
  input         io_decex_memOp_byte,
  input         io_decex_memOp_zext,
  input  [1:0]  io_decex_memOp_typ,
  input  [2:0]  io_decex_stackOp,
  input  [4:0]  io_decex_rsAddr_0,
  input  [4:0]  io_decex_rsAddr_1,
  input  [4:0]  io_decex_rsAddr_2,
  input  [4:0]  io_decex_rsAddr_3,
  input  [31:0] io_decex_rsData_0,
  input  [31:0] io_decex_rsData_1,
  input  [31:0] io_decex_rsData_2,
  input  [31:0] io_decex_rsData_3,
  input  [4:0]  io_decex_rdAddr_0,
  input  [4:0]  io_decex_rdAddr_1,
  input  [31:0] io_decex_immVal_0,
  input  [31:0] io_decex_immVal_1,
  input         io_decex_immOp_0,
  input         io_decex_immOp_1,
  input         io_decex_wrRd_0,
  input         io_decex_wrRd_1,
  input  [31:0] io_decex_callAddr,
  input         io_decex_call,
  input         io_decex_ret,
  input         io_decex_brcf,
  input         io_decex_trap,
  input         io_decex_xcall,
  input         io_decex_xret,
  input  [4:0]  io_decex_xsrc,
  input         io_decex_nonDelayed,
  input         io_decex_illOp,
  output [4:0]  io_exmem_rd_0_addr,
  output [31:0] io_exmem_rd_0_data,
  output        io_exmem_rd_0_valid,
  output [4:0]  io_exmem_rd_1_addr,
  output [31:0] io_exmem_rd_1_data,
  output        io_exmem_rd_1_valid,
  output        io_exmem_mem_load,
  output        io_exmem_mem_store,
  output        io_exmem_mem_hword,
  output        io_exmem_mem_byte,
  output        io_exmem_mem_zext,
  output [1:0]  io_exmem_mem_typ,
  output [31:0] io_exmem_mem_addr,
  output [31:0] io_exmem_mem_data,
  output        io_exmem_mem_call,
  output        io_exmem_mem_ret,
  output        io_exmem_mem_brcf,
  output        io_exmem_mem_trap,
  output        io_exmem_mem_xcall,
  output        io_exmem_mem_xret,
  output [4:0]  io_exmem_mem_xsrc,
  output        io_exmem_mem_illOp,
  output        io_exmem_mem_nonDelayed,
  output [29:0] io_exmem_base,
  output [29:0] io_exmem_relPc,
  output        io_exicache_doCallRet,
  output [31:0] io_exicache_callRetBase,
  output [31:0] io_exicache_callRetAddr,
  input  [29:0] io_feex_pc,
  input  [4:0]  io_exResult_0_addr,
  input  [31:0] io_exResult_0_data,
  input         io_exResult_0_valid,
  input  [4:0]  io_exResult_1_addr,
  input  [31:0] io_exResult_1_data,
  input         io_exResult_1_valid,
  input  [4:0]  io_memResult_0_addr,
  input  [31:0] io_memResult_0_data,
  input         io_memResult_0_valid,
  input  [4:0]  io_memResult_1_addr,
  input  [31:0] io_memResult_1_data,
  input         io_memResult_1_valid,
  output        io_exfe_doBranch,
  output [29:0] io_exfe_branchPc,
  output [2:0]  io_exsc_op,
  output [31:0] io_exsc_opData,
  output [31:0] io_exsc_opOff,
  input  [31:0] io_scex_stackTop,
  input  [31:0] io_scex_memTop
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
`endif // RANDOMIZE_REG_INIT
  reg [29:0] exReg_base; // @[Execute.scala 18:18]
  reg [29:0] exReg_relPc; // @[Execute.scala 18:18]
  reg [3:0] exReg_pred_0; // @[Execute.scala 18:18]
  reg [3:0] exReg_pred_1; // @[Execute.scala 18:18]
  reg [3:0] exReg_aluOp_0_func; // @[Execute.scala 18:18]
  reg  exReg_aluOp_0_isMul; // @[Execute.scala 18:18]
  reg  exReg_aluOp_0_isCmp; // @[Execute.scala 18:18]
  reg  exReg_aluOp_0_isPred; // @[Execute.scala 18:18]
  reg  exReg_aluOp_0_isBCpy; // @[Execute.scala 18:18]
  reg  exReg_aluOp_0_isMTS; // @[Execute.scala 18:18]
  reg  exReg_aluOp_0_isMFS; // @[Execute.scala 18:18]
  reg [3:0] exReg_aluOp_1_func; // @[Execute.scala 18:18]
  reg  exReg_aluOp_1_isCmp; // @[Execute.scala 18:18]
  reg  exReg_aluOp_1_isPred; // @[Execute.scala 18:18]
  reg  exReg_aluOp_1_isBCpy; // @[Execute.scala 18:18]
  reg  exReg_aluOp_1_isMTS; // @[Execute.scala 18:18]
  reg  exReg_aluOp_1_isMFS; // @[Execute.scala 18:18]
  reg [1:0] exReg_predOp_0_func; // @[Execute.scala 18:18]
  reg [2:0] exReg_predOp_0_dest; // @[Execute.scala 18:18]
  reg [3:0] exReg_predOp_0_s1Addr; // @[Execute.scala 18:18]
  reg [3:0] exReg_predOp_0_s2Addr; // @[Execute.scala 18:18]
  reg [1:0] exReg_predOp_1_func; // @[Execute.scala 18:18]
  reg [2:0] exReg_predOp_1_dest; // @[Execute.scala 18:18]
  reg [3:0] exReg_predOp_1_s1Addr; // @[Execute.scala 18:18]
  reg [3:0] exReg_predOp_1_s2Addr; // @[Execute.scala 18:18]
  reg  exReg_jmpOp_branch; // @[Execute.scala 18:18]
  reg [29:0] exReg_jmpOp_target; // @[Execute.scala 18:18]
  reg [31:0] exReg_jmpOp_reloc; // @[Execute.scala 18:18]
  reg  exReg_memOp_load; // @[Execute.scala 18:18]
  reg  exReg_memOp_store; // @[Execute.scala 18:18]
  reg  exReg_memOp_hword; // @[Execute.scala 18:18]
  reg  exReg_memOp_byte; // @[Execute.scala 18:18]
  reg  exReg_memOp_zext; // @[Execute.scala 18:18]
  reg [1:0] exReg_memOp_typ; // @[Execute.scala 18:18]
  reg [2:0] exReg_stackOp; // @[Execute.scala 18:18]
  reg [31:0] exReg_rsData_0; // @[Execute.scala 18:18]
  reg [31:0] exReg_rsData_1; // @[Execute.scala 18:18]
  reg [31:0] exReg_rsData_2; // @[Execute.scala 18:18]
  reg [31:0] exReg_rsData_3; // @[Execute.scala 18:18]
  reg [4:0] exReg_rdAddr_0; // @[Execute.scala 18:18]
  reg [4:0] exReg_rdAddr_1; // @[Execute.scala 18:18]
  reg [31:0] exReg_immVal_0; // @[Execute.scala 18:18]
  reg [31:0] exReg_immVal_1; // @[Execute.scala 18:18]
  reg  exReg_immOp_0; // @[Execute.scala 18:18]
  reg  exReg_wrRd_0; // @[Execute.scala 18:18]
  reg  exReg_wrRd_1; // @[Execute.scala 18:18]
  reg [31:0] exReg_callAddr; // @[Execute.scala 18:18]
  reg  exReg_call; // @[Execute.scala 18:18]
  reg  exReg_ret; // @[Execute.scala 18:18]
  reg  exReg_brcf; // @[Execute.scala 18:18]
  reg  exReg_trap; // @[Execute.scala 18:18]
  reg  exReg_xcall; // @[Execute.scala 18:18]
  reg  exReg_xret; // @[Execute.scala 18:18]
  reg [4:0] exReg_xsrc; // @[Execute.scala 18:18]
  reg  exReg_nonDelayed; // @[Execute.scala 18:18]
  reg  exReg_illOp; // @[Execute.scala 18:18]
  reg [2:0] fwReg_0; // @[Execute.scala 81:19]
  reg [2:0] fwReg_1; // @[Execute.scala 81:19]
  reg [2:0] fwReg_2; // @[Execute.scala 81:19]
  reg [2:0] fwReg_3; // @[Execute.scala 81:19]
  reg  fwSrcReg_0; // @[Execute.scala 82:22]
  reg  fwSrcReg_1; // @[Execute.scala 82:22]
  reg  fwSrcReg_2; // @[Execute.scala 82:22]
  reg  fwSrcReg_3; // @[Execute.scala 82:22]
  reg [31:0] memResultDataReg_0; // @[Execute.scala 83:29]
  reg [31:0] memResultDataReg_1; // @[Execute.scala 83:29]
  reg [31:0] exResultDataReg_0; // @[Execute.scala 84:29]
  reg [31:0] exResultDataReg_1; // @[Execute.scala 84:29]
  wire [2:0] _GEN_67 = io_decex_rsAddr_0 == io_memResult_0_addr & io_memResult_0_valid ? 3'h2 : 3'h0; // @[Execute.scala 92:82 Execute.scala 93:18 Execute.scala 89:14]
  wire  _T_6 = io_decex_rsAddr_0 == io_memResult_1_addr & io_memResult_1_valid; // @[Execute.scala 92:56]
  wire  _GEN_72 = io_decex_rsAddr_0 == io_exResult_0_addr & io_exResult_0_valid ? 1'h0 : _T_6; // @[Execute.scala 98:80 Execute.scala 100:21]
  wire  _GEN_74 = io_decex_rsAddr_0 == io_exResult_1_addr & io_exResult_1_valid | _GEN_72; // @[Execute.scala 98:80 Execute.scala 100:21]
  wire [2:0] _GEN_75 = io_decex_rsAddr_1 == io_memResult_0_addr & io_memResult_0_valid ? 3'h2 : 3'h0; // @[Execute.scala 92:82 Execute.scala 93:18 Execute.scala 89:14]
  wire  _T_14 = io_decex_rsAddr_1 == io_memResult_1_addr & io_memResult_1_valid; // @[Execute.scala 92:56]
  wire [2:0] _GEN_77 = io_decex_rsAddr_1 == io_memResult_1_addr & io_memResult_1_valid ? 3'h2 : _GEN_75; // @[Execute.scala 92:82 Execute.scala 93:18]
  wire  _GEN_80 = io_decex_rsAddr_1 == io_exResult_0_addr & io_exResult_0_valid ? 1'h0 : _T_14; // @[Execute.scala 98:80 Execute.scala 100:21]
  wire  _GEN_82 = io_decex_rsAddr_1 == io_exResult_1_addr & io_exResult_1_valid | _GEN_80; // @[Execute.scala 98:80 Execute.scala 100:21]
  wire [2:0] _GEN_83 = io_decex_rsAddr_2 == io_memResult_0_addr & io_memResult_0_valid ? 3'h2 : 3'h0; // @[Execute.scala 92:82 Execute.scala 93:18 Execute.scala 89:14]
  wire  _T_22 = io_decex_rsAddr_2 == io_memResult_1_addr & io_memResult_1_valid; // @[Execute.scala 92:56]
  wire  _GEN_88 = io_decex_rsAddr_2 == io_exResult_0_addr & io_exResult_0_valid ? 1'h0 : _T_22; // @[Execute.scala 98:80 Execute.scala 100:21]
  wire  _GEN_90 = io_decex_rsAddr_2 == io_exResult_1_addr & io_exResult_1_valid | _GEN_88; // @[Execute.scala 98:80 Execute.scala 100:21]
  wire [2:0] _GEN_91 = io_decex_rsAddr_3 == io_memResult_0_addr & io_memResult_0_valid ? 3'h2 : 3'h0; // @[Execute.scala 92:82 Execute.scala 93:18 Execute.scala 89:14]
  wire  _T_30 = io_decex_rsAddr_3 == io_memResult_1_addr & io_memResult_1_valid; // @[Execute.scala 92:56]
  wire [2:0] _GEN_93 = io_decex_rsAddr_3 == io_memResult_1_addr & io_memResult_1_valid ? 3'h2 : _GEN_91; // @[Execute.scala 92:82 Execute.scala 93:18]
  wire  _GEN_96 = io_decex_rsAddr_3 == io_exResult_0_addr & io_exResult_0_valid ? 1'h0 : _T_30; // @[Execute.scala 98:80 Execute.scala 100:21]
  wire  _GEN_98 = io_decex_rsAddr_3 == io_exResult_1_addr & io_exResult_1_valid | _GEN_96; // @[Execute.scala 98:80 Execute.scala 100:21]
  wire  _T_35 = ~io_ena; // @[Execute.scala 110:9]
  wire [31:0] _GEN_114 = fwSrcReg_0 ? memResultDataReg_1 : memResultDataReg_0; // @[Execute.scala 122:23 Execute.scala 122:23]
  wire [31:0] _T_38 = fwReg_0[1] ? _GEN_114 : exReg_rsData_0; // @[Execute.scala 122:23]
  wire [31:0] _GEN_116 = fwSrcReg_0 ? exResultDataReg_1 : exResultDataReg_0; // @[Execute.scala 121:19 Execute.scala 121:19]
  wire [31:0] op_0 = fwReg_0[0] ? _GEN_116 : _T_38; // @[Execute.scala 121:19]
  wire [31:0] _T_43 = fwReg_1[2] ? exReg_immVal_0 : exReg_rsData_1; // @[Execute.scala 127:29]
  wire [31:0] _GEN_118 = fwSrcReg_1 ? memResultDataReg_1 : memResultDataReg_0; // @[Execute.scala 126:25 Execute.scala 126:25]
  wire [31:0] _T_44 = fwReg_1[1] ? _GEN_118 : _T_43; // @[Execute.scala 126:25]
  wire [31:0] _GEN_120 = fwSrcReg_1 ? exResultDataReg_1 : exResultDataReg_0; // @[Execute.scala 125:21 Execute.scala 125:21]
  wire [31:0] op_1 = fwReg_1[0] ? _GEN_120 : _T_44; // @[Execute.scala 125:21]
  wire [31:0] _GEN_122 = fwSrcReg_2 ? memResultDataReg_1 : memResultDataReg_0; // @[Execute.scala 122:23 Execute.scala 122:23]
  wire [31:0] _T_48 = fwReg_2[1] ? _GEN_122 : exReg_rsData_2; // @[Execute.scala 122:23]
  wire [31:0] _GEN_124 = fwSrcReg_2 ? exResultDataReg_1 : exResultDataReg_0; // @[Execute.scala 121:19 Execute.scala 121:19]
  wire [31:0] op_2 = fwReg_2[0] ? _GEN_124 : _T_48; // @[Execute.scala 121:19]
  wire [31:0] _T_53 = fwReg_3[2] ? exReg_immVal_1 : exReg_rsData_3; // @[Execute.scala 127:29]
  wire [31:0] _GEN_126 = fwSrcReg_3 ? memResultDataReg_1 : memResultDataReg_0; // @[Execute.scala 126:25 Execute.scala 126:25]
  wire [31:0] _T_54 = fwReg_3[1] ? _GEN_126 : _T_53; // @[Execute.scala 126:25]
  wire [31:0] _GEN_128 = fwSrcReg_3 ? exResultDataReg_1 : exResultDataReg_0; // @[Execute.scala 125:21 Execute.scala 125:21]
  wire [31:0] op_3 = fwReg_3[0] ? _GEN_128 : _T_54; // @[Execute.scala 125:21]
  reg  predReg_1; // @[Execute.scala 132:20]
  reg  predReg_2; // @[Execute.scala 132:20]
  reg  predReg_3; // @[Execute.scala 132:20]
  reg  predReg_4; // @[Execute.scala 132:20]
  reg  predReg_5; // @[Execute.scala 132:20]
  reg  predReg_6; // @[Execute.scala 132:20]
  reg  predReg_7; // @[Execute.scala 132:20]
  wire  _GEN_130 = 3'h1 == exReg_pred_0[2:0] ? predReg_1 : 1'h1; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_131 = 3'h2 == exReg_pred_0[2:0] ? predReg_2 : _GEN_130; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_132 = 3'h3 == exReg_pred_0[2:0] ? predReg_3 : _GEN_131; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_133 = 3'h4 == exReg_pred_0[2:0] ? predReg_4 : _GEN_132; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_134 = 3'h5 == exReg_pred_0[2:0] ? predReg_5 : _GEN_133; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_135 = 3'h6 == exReg_pred_0[2:0] ? predReg_6 : _GEN_134; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_136 = 3'h7 == exReg_pred_0[2:0] ? predReg_7 : _GEN_135; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _T_58 = _GEN_136 ^ exReg_pred_0[3]; // @[Execute.scala 137:64]
  wire  doExecute_0 = io_flush ? 1'h0 : _T_58; // @[Execute.scala 136:24]
  wire  _GEN_138 = 3'h1 == exReg_pred_1[2:0] ? predReg_1 : 1'h1; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_139 = 3'h2 == exReg_pred_1[2:0] ? predReg_2 : _GEN_138; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_140 = 3'h3 == exReg_pred_1[2:0] ? predReg_3 : _GEN_139; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_141 = 3'h4 == exReg_pred_1[2:0] ? predReg_4 : _GEN_140; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_142 = 3'h5 == exReg_pred_1[2:0] ? predReg_5 : _GEN_141; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_143 = 3'h6 == exReg_pred_1[2:0] ? predReg_6 : _GEN_142; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _GEN_144 = 3'h7 == exReg_pred_1[2:0] ? predReg_7 : _GEN_143; // @[Execute.scala 137:64 Execute.scala 137:64]
  wire  _T_62 = _GEN_144 ^ exReg_pred_1[3]; // @[Execute.scala 137:64]
  wire  doExecute_1 = io_flush ? 1'h0 : _T_62; // @[Execute.scala 136:24]
  reg [31:0] retBaseReg; // @[Execute.scala 141:23]
  reg [31:0] retOffReg; // @[Execute.scala 142:22]
  reg  saveRetOff; // @[Execute.scala 143:23]
  reg  saveND; // @[Execute.scala 144:19]
  reg [31:0] excBaseReg; // @[Execute.scala 147:23]
  reg [31:0] excOffReg; // @[Execute.scala 148:22]
  reg [31:0] mulLoReg; // @[Execute.scala 153:21]
  reg [31:0] mulHiReg; // @[Execute.scala 154:21]
  reg [31:0] mulLLReg; // @[Execute.scala 157:24]
  reg [32:0] mulLHReg; // @[Execute.scala 158:24]
  reg [32:0] mulHLReg; // @[Execute.scala 159:24]
  reg [31:0] mulHHReg; // @[Execute.scala 160:24]
  reg  mulPipeReg; // @[Execute.scala 162:23]
  wire  _T_65 = exReg_aluOp_0_func == 4'h0; // @[Execute.scala 168:38]
  wire  hi = _T_65 & op_0[31]; // @[Execute.scala 170:23]
  wire [15:0] lo = op_0[31:16]; // @[Execute.scala 171:25]
  wire [16:0] _T_68 = {hi,lo}; // @[Execute.scala 171:55]
  wire  hi_1 = _T_65 & op_1[31]; // @[Execute.scala 173:23]
  wire [15:0] lo_1 = op_1[31:16]; // @[Execute.scala 174:25]
  wire [16:0] _T_72 = {hi_1,lo_1}; // @[Execute.scala 174:55]
  wire [31:0] _T_74 = op_0[15:0] * op_1[15:0]; // @[Execute.scala 177:22]
  wire [16:0] _T_75 = {1'b0,$signed(op_0[15:0])}; // @[Execute.scala 178:22]
  wire [33:0] _T_76 = $signed(_T_72) * $signed(_T_75); // @[Execute.scala 178:22]
  wire [32:0] _T_78 = _T_76[32:0]; // @[Execute.scala 178:22]
  wire [16:0] _T_79 = {1'b0,$signed(op_1[15:0])}; // @[Execute.scala 179:22]
  wire [33:0] _T_80 = $signed(_T_68) * $signed(_T_79); // @[Execute.scala 179:22]
  wire [32:0] _T_82 = _T_80[32:0]; // @[Execute.scala 179:22]
  wire [33:0] _T_84 = $signed(_T_68) * $signed(_T_72); // @[Execute.scala 180:31]
  wire [63:0] _T_86 = {mulHHReg,mulLLReg}; // @[Execute.scala 182:46]
  wire [48:0] _T_88 = {mulHLReg,16'h0}; // @[Execute.scala 183:69]
  wire [63:0] _GEN_423 = {{15{_T_88[48]}},_T_88}; // @[Execute.scala 183:22]
  wire [63:0] _T_91 = $signed(_T_86) + $signed(_GEN_423); // @[Execute.scala 183:22]
  wire [48:0] _T_93 = {mulLHReg,16'h0}; // @[Execute.scala 184:69]
  wire [63:0] _GEN_424 = {{15{_T_93[48]}},_T_93}; // @[Execute.scala 184:22]
  wire [63:0] _T_96 = $signed(_T_91) + $signed(_GEN_424); // @[Execute.scala 184:22]
  wire [31:0] _GEN_145 = mulPipeReg ? _T_96[63:32] : mulHiReg; // @[Execute.scala 186:22 Execute.scala 187:16 Execute.scala 154:21]
  wire [31:0] _GEN_146 = mulPipeReg ? _T_96[31:0] : mulLoReg; // @[Execute.scala 186:22 Execute.scala 188:16 Execute.scala 153:21]
  wire [33:0] _GEN_151 = io_ena ? _T_84 : {{2'd0}, mulHHReg}; // @[Execute.scala 165:16 Execute.scala 180:14 Execute.scala 160:24]
  wire [31:0] _GEN_152 = io_ena ? _GEN_145 : mulHiReg; // @[Execute.scala 165:16 Execute.scala 154:21]
  wire [31:0] _GEN_153 = io_ena ? _GEN_146 : mulLoReg; // @[Execute.scala 165:16 Execute.scala 153:21]
  wire [2:0] _GEN_154 = ~io_brflush & doExecute_0 ? exReg_stackOp : 3'h0; // @[Execute.scala 198:37 Execute.scala 199:16 Execute.scala 193:14]
  wire  _T_103 = exReg_aluOp_0_func == 4'hc; // @[Execute.scala 30:41]
  wire [1:0] _T_105 = exReg_aluOp_0_func == 4'hd ? 2'h2 : {{1'd0}, _T_103}; // @[Execute.scala 29:31]
  wire [34:0] _GEN_425 = {{3'd0}, op_0}; // @[Execute.scala 29:25]
  wire [34:0] _T_106 = _GEN_425 << _T_105; // @[Execute.scala 29:25]
  wire [34:0] _GEN_426 = {{3'd0}, op_1}; // @[Execute.scala 32:25]
  wire [34:0] _T_108 = _T_106 + _GEN_426; // @[Execute.scala 32:25]
  wire  _T_112 = exReg_aluOp_0_func == 4'h5 & op_0[31]; // @[Execute.scala 35:19]
  wire  _T_114 = 4'h0 == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire  _T_115 = 4'h1 == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire [31:0] _T_117 = op_0 - op_1; // @[Execute.scala 40:39]
  wire  _T_118 = 4'h2 == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire [31:0] _T_119 = op_0 ^ op_1; // @[Execute.scala 41:40]
  wire  _T_120 = 4'h3 == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire [62:0] _GEN_427 = {{31'd0}, op_0}; // @[Execute.scala 42:40]
  wire [62:0] _T_121 = _GEN_427 << op_1[4:0]; // @[Execute.scala 42:40]
  wire  _T_123 = 4'h4 == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire  _T_124 = 4'h5 == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire  _T_125 = 4'h4 == exReg_aluOp_0_func | 4'h5 == exReg_aluOp_0_func; // @[Conditional.scala 37:55]
  wire [32:0] _T_126 = {_T_112,op_0}; // @[Execute.scala 43:47]
  wire [32:0] _T_128 = $signed(_T_126) >>> op_1[4:0]; // @[Execute.scala 43:64]
  wire  _T_129 = 4'h6 == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire [31:0] _T_130 = op_0 | op_1; // @[Execute.scala 44:40]
  wire  _T_131 = 4'h7 == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire [31:0] _T_132 = op_0 & op_1; // @[Execute.scala 45:40]
  wire  _T_133 = 4'hb == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire [31:0] _T_135 = ~_T_130; // @[Execute.scala 46:36]
  wire [34:0] _GEN_157 = _T_133 ? {{3'd0}, _T_135} : _T_108; // @[Conditional.scala 39:67 Execute.scala 46:32]
  wire [34:0] _GEN_158 = _T_131 ? {{3'd0}, _T_132} : _GEN_157; // @[Conditional.scala 39:67 Execute.scala 45:32]
  wire [34:0] _GEN_159 = _T_129 ? {{3'd0}, _T_130} : _GEN_158; // @[Conditional.scala 39:67 Execute.scala 44:32]
  wire [34:0] _GEN_160 = _T_125 ? {{2'd0}, _T_128} : _GEN_159; // @[Conditional.scala 39:67 Execute.scala 43:38]
  wire [34:0] _GEN_161 = _T_120 ? {{3'd0}, _T_121[31:0]} : _GEN_160; // @[Conditional.scala 39:67 Execute.scala 42:32]
  wire [34:0] _GEN_162 = _T_118 ? {{3'd0}, _T_119} : _GEN_161; // @[Conditional.scala 39:67 Execute.scala 41:32]
  wire [34:0] _GEN_163 = _T_115 ? {{3'd0}, _T_117} : _GEN_162; // @[Conditional.scala 39:67 Execute.scala 40:32]
  wire [34:0] _GEN_164 = _T_114 ? _T_108 : _GEN_163; // @[Conditional.scala 40:58 Execute.scala 39:32]
  wire [31:0] _T_138 = fwReg_0[0] ? _GEN_116 : _T_38; // @[Execute.scala 54:20]
  wire [31:0] _T_139 = fwReg_1[0] ? _GEN_120 : _T_44; // @[Execute.scala 55:20]
  wire [31:0] _T_141 = 32'h1 << op_1[4:0]; // @[Execute.scala 56:26]
  wire  _T_142 = op_0 == op_1; // @[Execute.scala 59:18]
  wire  _T_143 = $signed(_T_138) < $signed(_T_139); // @[Execute.scala 60:19]
  wire  _T_144 = op_0 < op_1; // @[Execute.scala 61:19]
  wire  _T_145 = ~_T_142; // @[Execute.scala 64:21]
  wire  _T_146 = _T_143 | _T_142; // @[Execute.scala 66:24]
  wire  _T_147 = _T_144 | _T_142; // @[Execute.scala 68:25]
  wire [31:0] _T_148 = op_0 & _T_141; // @[Execute.scala 69:26]
  wire  _T_149 = _T_148 != 32'h0; // @[Execute.scala 69:36]
  wire  _T_153 = _T_115 ? _T_145 : _T_114 & _T_142; // @[Mux.scala 80:57]
  wire  _T_155 = _T_118 ? _T_143 : _T_153; // @[Mux.scala 80:57]
  wire  _T_157 = _T_120 ? _T_146 : _T_155; // @[Mux.scala 80:57]
  wire  _T_159 = _T_123 ? _T_144 : _T_157; // @[Mux.scala 80:57]
  wire  _T_161 = _T_124 ? _T_147 : _T_159; // @[Mux.scala 80:57]
  wire  _T_163 = _T_129 ? _T_149 : _T_161; // @[Mux.scala 80:57]
  wire  _GEN_166 = 3'h1 == exReg_aluOp_0_func[2:0] ? predReg_1 : 1'h1; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_167 = 3'h2 == exReg_aluOp_0_func[2:0] ? predReg_2 : _GEN_166; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_168 = 3'h3 == exReg_aluOp_0_func[2:0] ? predReg_3 : _GEN_167; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_169 = 3'h4 == exReg_aluOp_0_func[2:0] ? predReg_4 : _GEN_168; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_170 = 3'h5 == exReg_aluOp_0_func[2:0] ? predReg_5 : _GEN_169; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_171 = 3'h6 == exReg_aluOp_0_func[2:0] ? predReg_6 : _GEN_170; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_172 = 3'h7 == exReg_aluOp_0_func[2:0] ? predReg_7 : _GEN_171; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _T_166 = _GEN_172 ^ exReg_aluOp_0_func[3]; // @[Execute.scala 208:63]
  wire [31:0] _T_167 = {31'h0,_T_166}; // @[Execute.scala 209:45]
  wire [62:0] _GEN_428 = {{31'd0}, _T_167}; // @[Execute.scala 209:56]
  wire [62:0] _T_169 = _GEN_428 << op_1[4:0]; // @[Execute.scala 209:56]
  wire [62:0] _T_172 = 63'h1 << op_1[4:0]; // @[Execute.scala 210:60]
  wire [31:0] _T_174 = ~_T_172[31:0]; // @[Execute.scala 210:30]
  wire [31:0] _T_175 = op_0 & _T_174; // @[Execute.scala 210:28]
  wire [31:0] _T_176 = _T_175 | _T_169[31:0]; // @[Execute.scala 211:31]
  wire  _GEN_174 = 3'h1 == exReg_predOp_0_s1Addr[2:0] ? predReg_1 : 1'h1; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_175 = 3'h2 == exReg_predOp_0_s1Addr[2:0] ? predReg_2 : _GEN_174; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_176 = 3'h3 == exReg_predOp_0_s1Addr[2:0] ? predReg_3 : _GEN_175; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_177 = 3'h4 == exReg_predOp_0_s1Addr[2:0] ? predReg_4 : _GEN_176; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_178 = 3'h5 == exReg_predOp_0_s1Addr[2:0] ? predReg_5 : _GEN_177; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_179 = 3'h6 == exReg_predOp_0_s1Addr[2:0] ? predReg_6 : _GEN_178; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_180 = 3'h7 == exReg_predOp_0_s1Addr[2:0] ? predReg_7 : _GEN_179; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _T_179 = _GEN_180 ^ exReg_predOp_0_s1Addr[3]; // @[Execute.scala 214:62]
  wire  _GEN_182 = 3'h1 == exReg_predOp_0_s2Addr[2:0] ? predReg_1 : 1'h1; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_183 = 3'h2 == exReg_predOp_0_s2Addr[2:0] ? predReg_2 : _GEN_182; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_184 = 3'h3 == exReg_predOp_0_s2Addr[2:0] ? predReg_3 : _GEN_183; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_185 = 3'h4 == exReg_predOp_0_s2Addr[2:0] ? predReg_4 : _GEN_184; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_186 = 3'h5 == exReg_predOp_0_s2Addr[2:0] ? predReg_5 : _GEN_185; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_187 = 3'h6 == exReg_predOp_0_s2Addr[2:0] ? predReg_6 : _GEN_186; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_188 = 3'h7 == exReg_predOp_0_s2Addr[2:0] ? predReg_7 : _GEN_187; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _T_182 = _GEN_188 ^ exReg_predOp_0_s2Addr[3]; // @[Execute.scala 215:62]
  wire  _T_183 = _T_179 | _T_182; // @[Execute.scala 74:22]
  wire  _T_184 = _T_179 & _T_182; // @[Execute.scala 75:23]
  wire  _T_185 = _T_179 ^ _T_182; // @[Execute.scala 76:23]
  wire  _T_187 = ~_T_183; // @[Execute.scala 77:19]
  wire  _T_189 = 2'h1 == exReg_predOp_0_func ? _T_184 : _T_183; // @[Mux.scala 80:57]
  wire  _T_191 = 2'h2 == exReg_predOp_0_func ? _T_185 : _T_189; // @[Mux.scala 80:57]
  wire  _T_193 = 2'h3 == exReg_predOp_0_func ? _T_187 : _T_191; // @[Mux.scala 80:57]
  wire  _T_196 = exReg_aluOp_0_isCmp ? _T_163 : _T_193; // @[Execute.scala 219:43]
  wire  _GEN_190 = 3'h1 == exReg_predOp_0_dest ? _T_196 : predReg_1; // @[Execute.scala 219:37 Execute.scala 219:37 Execute.scala 132:20]
  wire  _GEN_191 = 3'h2 == exReg_predOp_0_dest ? _T_196 : predReg_2; // @[Execute.scala 219:37 Execute.scala 219:37 Execute.scala 132:20]
  wire  _GEN_192 = 3'h3 == exReg_predOp_0_dest ? _T_196 : predReg_3; // @[Execute.scala 219:37 Execute.scala 219:37 Execute.scala 132:20]
  wire  _GEN_193 = 3'h4 == exReg_predOp_0_dest ? _T_196 : predReg_4; // @[Execute.scala 219:37 Execute.scala 219:37 Execute.scala 132:20]
  wire  _GEN_194 = 3'h5 == exReg_predOp_0_dest ? _T_196 : predReg_5; // @[Execute.scala 219:37 Execute.scala 219:37 Execute.scala 132:20]
  wire  _GEN_195 = 3'h6 == exReg_predOp_0_dest ? _T_196 : predReg_6; // @[Execute.scala 219:37 Execute.scala 219:37 Execute.scala 132:20]
  wire  _GEN_196 = 3'h7 == exReg_predOp_0_dest ? _T_196 : predReg_7; // @[Execute.scala 219:37 Execute.scala 219:37 Execute.scala 132:20]
  wire  _GEN_198 = (exReg_aluOp_0_isCmp | exReg_aluOp_0_isPred) & doExecute_0 ? _GEN_190 : predReg_1; // @[Execute.scala 218:75 Execute.scala 132:20]
  wire  _GEN_199 = (exReg_aluOp_0_isCmp | exReg_aluOp_0_isPred) & doExecute_0 ? _GEN_191 : predReg_2; // @[Execute.scala 218:75 Execute.scala 132:20]
  wire  _GEN_200 = (exReg_aluOp_0_isCmp | exReg_aluOp_0_isPred) & doExecute_0 ? _GEN_192 : predReg_3; // @[Execute.scala 218:75 Execute.scala 132:20]
  wire  _GEN_201 = (exReg_aluOp_0_isCmp | exReg_aluOp_0_isPred) & doExecute_0 ? _GEN_193 : predReg_4; // @[Execute.scala 218:75 Execute.scala 132:20]
  wire  _GEN_202 = (exReg_aluOp_0_isCmp | exReg_aluOp_0_isPred) & doExecute_0 ? _GEN_194 : predReg_5; // @[Execute.scala 218:75 Execute.scala 132:20]
  wire  _GEN_203 = (exReg_aluOp_0_isCmp | exReg_aluOp_0_isPred) & doExecute_0 ? _GEN_195 : predReg_6; // @[Execute.scala 218:75 Execute.scala 132:20]
  wire  _GEN_204 = (exReg_aluOp_0_isCmp | exReg_aluOp_0_isPred) & doExecute_0 ? _GEN_196 : predReg_7; // @[Execute.scala 218:75 Execute.scala 132:20]
  wire  _T_212 = 4'h8 == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire  _T_213 = 4'h9 == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire  _T_214 = 4'ha == exReg_aluOp_0_func; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_205 = _T_214 ? op_0 : excOffReg; // @[Conditional.scala 39:67 Execute.scala 257:21 Execute.scala 148:22]
  wire [31:0] _GEN_206 = _T_213 ? op_0 : excBaseReg; // @[Conditional.scala 39:67 Execute.scala 254:22 Execute.scala 147:23]
  wire [31:0] _GEN_207 = _T_213 ? excOffReg : _GEN_205; // @[Conditional.scala 39:67 Execute.scala 148:22]
  wire [31:0] _GEN_208 = _T_212 ? op_0 : retOffReg; // @[Conditional.scala 39:67 Execute.scala 251:21 Execute.scala 142:22]
  wire [31:0] _GEN_209 = _T_212 ? excBaseReg : _GEN_206; // @[Conditional.scala 39:67 Execute.scala 147:23]
  wire [31:0] _GEN_210 = _T_212 ? excOffReg : _GEN_207; // @[Conditional.scala 39:67 Execute.scala 148:22]
  wire [31:0] _GEN_211 = _T_131 ? op_0 : retBaseReg; // @[Conditional.scala 39:67 Execute.scala 248:22 Execute.scala 141:23]
  wire [31:0] _GEN_212 = _T_131 ? retOffReg : _GEN_208; // @[Conditional.scala 39:67 Execute.scala 142:22]
  wire [31:0] _GEN_213 = _T_131 ? excBaseReg : _GEN_209; // @[Conditional.scala 39:67 Execute.scala 147:23]
  wire [31:0] _GEN_214 = _T_131 ? excOffReg : _GEN_210; // @[Conditional.scala 39:67 Execute.scala 148:22]
  wire [2:0] _GEN_215 = _T_124 ? 3'h2 : _GEN_154; // @[Conditional.scala 39:67 Execute.scala 245:22]
  wire [31:0] _GEN_216 = _T_124 ? retBaseReg : _GEN_211; // @[Conditional.scala 39:67 Execute.scala 141:23]
  wire [31:0] _GEN_217 = _T_124 ? retOffReg : _GEN_212; // @[Conditional.scala 39:67 Execute.scala 142:22]
  wire [31:0] _GEN_218 = _T_124 ? excBaseReg : _GEN_213; // @[Conditional.scala 39:67 Execute.scala 147:23]
  wire [31:0] _GEN_219 = _T_124 ? excOffReg : _GEN_214; // @[Conditional.scala 39:67 Execute.scala 148:22]
  wire [2:0] _GEN_220 = _T_129 ? 3'h1 : _GEN_215; // @[Conditional.scala 39:67 Execute.scala 242:22]
  wire [31:0] _GEN_221 = _T_129 ? retBaseReg : _GEN_216; // @[Conditional.scala 39:67 Execute.scala 141:23]
  wire [31:0] _GEN_222 = _T_129 ? retOffReg : _GEN_217; // @[Conditional.scala 39:67 Execute.scala 142:22]
  wire [31:0] _GEN_223 = _T_129 ? excBaseReg : _GEN_218; // @[Conditional.scala 39:67 Execute.scala 147:23]
  wire [31:0] _GEN_224 = _T_129 ? excOffReg : _GEN_219; // @[Conditional.scala 39:67 Execute.scala 148:22]
  wire [31:0] _GEN_225 = _T_120 ? op_0 : _GEN_152; // @[Conditional.scala 39:67 Execute.scala 239:20]
  wire [2:0] _GEN_226 = _T_120 ? _GEN_154 : _GEN_220; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_227 = _T_120 ? retBaseReg : _GEN_221; // @[Conditional.scala 39:67 Execute.scala 141:23]
  wire [31:0] _GEN_228 = _T_120 ? retOffReg : _GEN_222; // @[Conditional.scala 39:67 Execute.scala 142:22]
  wire [31:0] _GEN_229 = _T_120 ? excBaseReg : _GEN_223; // @[Conditional.scala 39:67 Execute.scala 147:23]
  wire [31:0] _GEN_230 = _T_120 ? excOffReg : _GEN_224; // @[Conditional.scala 39:67 Execute.scala 148:22]
  wire [31:0] _GEN_231 = _T_118 ? op_0 : _GEN_153; // @[Conditional.scala 39:67 Execute.scala 236:20]
  wire [31:0] _GEN_232 = _T_118 ? _GEN_152 : _GEN_225; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_233 = _T_118 ? _GEN_154 : _GEN_226; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_234 = _T_118 ? retBaseReg : _GEN_227; // @[Conditional.scala 39:67 Execute.scala 141:23]
  wire [31:0] _GEN_235 = _T_118 ? retOffReg : _GEN_228; // @[Conditional.scala 39:67 Execute.scala 142:22]
  wire [31:0] _GEN_236 = _T_118 ? excBaseReg : _GEN_229; // @[Conditional.scala 39:67 Execute.scala 147:23]
  wire [31:0] _GEN_237 = _T_118 ? excOffReg : _GEN_230; // @[Conditional.scala 39:67 Execute.scala 148:22]
  wire  _GEN_239 = _T_114 ? op_0[1] : _GEN_198; // @[Conditional.scala 40:58 Execute.scala 230:24]
  wire  _GEN_240 = _T_114 ? op_0[2] : _GEN_199; // @[Conditional.scala 40:58 Execute.scala 230:24]
  wire  _GEN_241 = _T_114 ? op_0[3] : _GEN_200; // @[Conditional.scala 40:58 Execute.scala 230:24]
  wire  _GEN_242 = _T_114 ? op_0[4] : _GEN_201; // @[Conditional.scala 40:58 Execute.scala 230:24]
  wire  _GEN_243 = _T_114 ? op_0[5] : _GEN_202; // @[Conditional.scala 40:58 Execute.scala 230:24]
  wire  _GEN_244 = _T_114 ? op_0[6] : _GEN_203; // @[Conditional.scala 40:58 Execute.scala 230:24]
  wire  _GEN_245 = _T_114 ? op_0[7] : _GEN_204; // @[Conditional.scala 40:58 Execute.scala 230:24]
  wire [31:0] _GEN_246 = _T_114 ? _GEN_153 : _GEN_231; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_247 = _T_114 ? _GEN_152 : _GEN_232; // @[Conditional.scala 40:58]
  wire [2:0] _GEN_248 = _T_114 ? _GEN_154 : _GEN_233; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_249 = _T_114 ? retBaseReg : _GEN_234; // @[Conditional.scala 40:58 Execute.scala 141:23]
  wire [31:0] _GEN_250 = _T_114 ? retOffReg : _GEN_235; // @[Conditional.scala 40:58 Execute.scala 142:22]
  wire [31:0] _GEN_251 = _T_114 ? excBaseReg : _GEN_236; // @[Conditional.scala 40:58 Execute.scala 147:23]
  wire [31:0] _GEN_252 = _T_114 ? excOffReg : _GEN_237; // @[Conditional.scala 40:58 Execute.scala 148:22]
  wire [31:0] _GEN_253 = exReg_aluOp_0_isMTS & doExecute_0 ? op_0 : 32'h0; // @[Execute.scala 224:48 Execute.scala 225:22 Execute.scala 194:18]
  wire  _GEN_255 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_239 : _GEN_198; // @[Execute.scala 224:48]
  wire  _GEN_256 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_240 : _GEN_199; // @[Execute.scala 224:48]
  wire  _GEN_257 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_241 : _GEN_200; // @[Execute.scala 224:48]
  wire  _GEN_258 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_242 : _GEN_201; // @[Execute.scala 224:48]
  wire  _GEN_259 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_243 : _GEN_202; // @[Execute.scala 224:48]
  wire  _GEN_260 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_244 : _GEN_203; // @[Execute.scala 224:48]
  wire  _GEN_261 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_245 : _GEN_204; // @[Execute.scala 224:48]
  wire [31:0] _GEN_262 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_246 : _GEN_153; // @[Execute.scala 224:48]
  wire [31:0] _GEN_263 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_247 : _GEN_152; // @[Execute.scala 224:48]
  wire [2:0] _GEN_264 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_248 : _GEN_154; // @[Execute.scala 224:48]
  wire [31:0] _GEN_265 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_249 : retBaseReg; // @[Execute.scala 224:48 Execute.scala 141:23]
  wire [31:0] _GEN_266 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_250 : retOffReg; // @[Execute.scala 224:48 Execute.scala 142:22]
  wire [31:0] _GEN_267 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_251 : excBaseReg; // @[Execute.scala 224:48 Execute.scala 147:23]
  wire [31:0] _GEN_268 = exReg_aluOp_0_isMTS & doExecute_0 ? _GEN_252 : excOffReg; // @[Execute.scala 224:48 Execute.scala 148:22]
  wire [31:0] _T_216 = {24'h0,predReg_7,predReg_6,predReg_5,predReg_4,predReg_3,predReg_2,predReg_1,1'h1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_269 = _T_214 ? excOffReg : 32'h0; // @[Conditional.scala 39:67 Execute.scala 289:19 Execute.scala 262:15]
  wire [31:0] _GEN_270 = _T_213 ? excBaseReg : _GEN_269; // @[Conditional.scala 39:67 Execute.scala 286:19]
  wire [31:0] _GEN_271 = _T_212 ? retOffReg : _GEN_270; // @[Conditional.scala 39:67 Execute.scala 283:19]
  wire [31:0] _GEN_272 = _T_131 ? retBaseReg : _GEN_271; // @[Conditional.scala 39:67 Execute.scala 280:19]
  wire [31:0] _GEN_273 = _T_124 ? io_scex_memTop : _GEN_272; // @[Conditional.scala 39:67 Execute.scala 277:19]
  wire [31:0] _GEN_274 = _T_129 ? io_scex_stackTop : _GEN_273; // @[Conditional.scala 39:67 Execute.scala 274:19]
  wire [31:0] _GEN_275 = _T_120 ? mulHiReg : _GEN_274; // @[Conditional.scala 39:67 Execute.scala 271:19]
  wire [31:0] _GEN_276 = _T_118 ? mulLoReg : _GEN_275; // @[Conditional.scala 39:67 Execute.scala 268:19]
  wire [31:0] _GEN_277 = _T_114 ? _T_216 : _GEN_276; // @[Conditional.scala 40:58 Execute.scala 265:19]
  wire [31:0] _T_226 = exReg_aluOp_0_isBCpy ? _T_176 : _GEN_164[31:0]; // @[Execute.scala 297:35]
  wire  _T_229 = exReg_aluOp_1_func == 4'hc; // @[Execute.scala 30:41]
  wire [1:0] _T_231 = exReg_aluOp_1_func == 4'hd ? 2'h2 : {{1'd0}, _T_229}; // @[Execute.scala 29:31]
  wire [34:0] _GEN_429 = {{3'd0}, op_2}; // @[Execute.scala 29:25]
  wire [34:0] _T_232 = _GEN_429 << _T_231; // @[Execute.scala 29:25]
  wire [34:0] _GEN_430 = {{3'd0}, op_3}; // @[Execute.scala 32:25]
  wire [34:0] _T_234 = _T_232 + _GEN_430; // @[Execute.scala 32:25]
  wire  _T_238 = exReg_aluOp_1_func == 4'h5 & op_2[31]; // @[Execute.scala 35:19]
  wire  _T_240 = 4'h0 == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire  _T_241 = 4'h1 == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire [31:0] _T_243 = op_2 - op_3; // @[Execute.scala 40:39]
  wire  _T_244 = 4'h2 == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire [31:0] _T_245 = op_2 ^ op_3; // @[Execute.scala 41:40]
  wire  _T_246 = 4'h3 == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire [62:0] _GEN_431 = {{31'd0}, op_2}; // @[Execute.scala 42:40]
  wire [62:0] _T_247 = _GEN_431 << op_3[4:0]; // @[Execute.scala 42:40]
  wire  _T_249 = 4'h4 == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire  _T_250 = 4'h5 == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire  _T_251 = 4'h4 == exReg_aluOp_1_func | 4'h5 == exReg_aluOp_1_func; // @[Conditional.scala 37:55]
  wire [32:0] _T_252 = {_T_238,op_2}; // @[Execute.scala 43:47]
  wire [32:0] _T_254 = $signed(_T_252) >>> op_3[4:0]; // @[Execute.scala 43:64]
  wire  _T_255 = 4'h6 == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire [31:0] _T_256 = op_2 | op_3; // @[Execute.scala 44:40]
  wire  _T_257 = 4'h7 == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire [31:0] _T_258 = op_2 & op_3; // @[Execute.scala 45:40]
  wire  _T_259 = 4'hb == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire [31:0] _T_261 = ~_T_256; // @[Execute.scala 46:36]
  wire [34:0] _GEN_280 = _T_259 ? {{3'd0}, _T_261} : _T_234; // @[Conditional.scala 39:67 Execute.scala 46:32]
  wire [34:0] _GEN_281 = _T_257 ? {{3'd0}, _T_258} : _GEN_280; // @[Conditional.scala 39:67 Execute.scala 45:32]
  wire [34:0] _GEN_282 = _T_255 ? {{3'd0}, _T_256} : _GEN_281; // @[Conditional.scala 39:67 Execute.scala 44:32]
  wire [34:0] _GEN_283 = _T_251 ? {{2'd0}, _T_254} : _GEN_282; // @[Conditional.scala 39:67 Execute.scala 43:38]
  wire [34:0] _GEN_284 = _T_246 ? {{3'd0}, _T_247[31:0]} : _GEN_283; // @[Conditional.scala 39:67 Execute.scala 42:32]
  wire [34:0] _GEN_285 = _T_244 ? {{3'd0}, _T_245} : _GEN_284; // @[Conditional.scala 39:67 Execute.scala 41:32]
  wire [34:0] _GEN_286 = _T_241 ? {{3'd0}, _T_243} : _GEN_285; // @[Conditional.scala 39:67 Execute.scala 40:32]
  wire [34:0] _GEN_287 = _T_240 ? _T_234 : _GEN_286; // @[Conditional.scala 40:58 Execute.scala 39:32]
  wire [31:0] _T_264 = fwReg_2[0] ? _GEN_124 : _T_48; // @[Execute.scala 54:20]
  wire [31:0] _T_265 = fwReg_3[0] ? _GEN_128 : _T_54; // @[Execute.scala 55:20]
  wire [31:0] _T_267 = 32'h1 << op_3[4:0]; // @[Execute.scala 56:26]
  wire  _T_268 = op_2 == op_3; // @[Execute.scala 59:18]
  wire  _T_269 = $signed(_T_264) < $signed(_T_265); // @[Execute.scala 60:19]
  wire  _T_270 = op_2 < op_3; // @[Execute.scala 61:19]
  wire  _T_271 = ~_T_268; // @[Execute.scala 64:21]
  wire  _T_272 = _T_269 | _T_268; // @[Execute.scala 66:24]
  wire  _T_273 = _T_270 | _T_268; // @[Execute.scala 68:25]
  wire [31:0] _T_274 = op_2 & _T_267; // @[Execute.scala 69:26]
  wire  _T_275 = _T_274 != 32'h0; // @[Execute.scala 69:36]
  wire  _T_279 = _T_241 ? _T_271 : _T_240 & _T_268; // @[Mux.scala 80:57]
  wire  _T_281 = _T_244 ? _T_269 : _T_279; // @[Mux.scala 80:57]
  wire  _T_283 = _T_246 ? _T_272 : _T_281; // @[Mux.scala 80:57]
  wire  _T_285 = _T_249 ? _T_270 : _T_283; // @[Mux.scala 80:57]
  wire  _T_287 = _T_250 ? _T_273 : _T_285; // @[Mux.scala 80:57]
  wire  _T_289 = _T_255 ? _T_275 : _T_287; // @[Mux.scala 80:57]
  wire  _GEN_289 = 3'h1 == exReg_aluOp_1_func[2:0] ? predReg_1 : 1'h1; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_290 = 3'h2 == exReg_aluOp_1_func[2:0] ? predReg_2 : _GEN_289; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_291 = 3'h3 == exReg_aluOp_1_func[2:0] ? predReg_3 : _GEN_290; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_292 = 3'h4 == exReg_aluOp_1_func[2:0] ? predReg_4 : _GEN_291; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_293 = 3'h5 == exReg_aluOp_1_func[2:0] ? predReg_5 : _GEN_292; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_294 = 3'h6 == exReg_aluOp_1_func[2:0] ? predReg_6 : _GEN_293; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _GEN_295 = 3'h7 == exReg_aluOp_1_func[2:0] ? predReg_7 : _GEN_294; // @[Execute.scala 208:63 Execute.scala 208:63]
  wire  _T_292 = _GEN_295 ^ exReg_aluOp_1_func[3]; // @[Execute.scala 208:63]
  wire [31:0] _T_293 = {31'h0,_T_292}; // @[Execute.scala 209:45]
  wire [62:0] _GEN_432 = {{31'd0}, _T_293}; // @[Execute.scala 209:56]
  wire [62:0] _T_295 = _GEN_432 << op_3[4:0]; // @[Execute.scala 209:56]
  wire [62:0] _T_298 = 63'h1 << op_3[4:0]; // @[Execute.scala 210:60]
  wire [31:0] _T_300 = ~_T_298[31:0]; // @[Execute.scala 210:30]
  wire [31:0] _T_301 = op_2 & _T_300; // @[Execute.scala 210:28]
  wire [31:0] _T_302 = _T_301 | _T_295[31:0]; // @[Execute.scala 211:31]
  wire  _GEN_297 = 3'h1 == exReg_predOp_1_s1Addr[2:0] ? predReg_1 : 1'h1; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_298 = 3'h2 == exReg_predOp_1_s1Addr[2:0] ? predReg_2 : _GEN_297; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_299 = 3'h3 == exReg_predOp_1_s1Addr[2:0] ? predReg_3 : _GEN_298; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_300 = 3'h4 == exReg_predOp_1_s1Addr[2:0] ? predReg_4 : _GEN_299; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_301 = 3'h5 == exReg_predOp_1_s1Addr[2:0] ? predReg_5 : _GEN_300; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_302 = 3'h6 == exReg_predOp_1_s1Addr[2:0] ? predReg_6 : _GEN_301; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _GEN_303 = 3'h7 == exReg_predOp_1_s1Addr[2:0] ? predReg_7 : _GEN_302; // @[Execute.scala 214:62 Execute.scala 214:62]
  wire  _T_305 = _GEN_303 ^ exReg_predOp_1_s1Addr[3]; // @[Execute.scala 214:62]
  wire  _GEN_305 = 3'h1 == exReg_predOp_1_s2Addr[2:0] ? predReg_1 : 1'h1; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_306 = 3'h2 == exReg_predOp_1_s2Addr[2:0] ? predReg_2 : _GEN_305; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_307 = 3'h3 == exReg_predOp_1_s2Addr[2:0] ? predReg_3 : _GEN_306; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_308 = 3'h4 == exReg_predOp_1_s2Addr[2:0] ? predReg_4 : _GEN_307; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_309 = 3'h5 == exReg_predOp_1_s2Addr[2:0] ? predReg_5 : _GEN_308; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_310 = 3'h6 == exReg_predOp_1_s2Addr[2:0] ? predReg_6 : _GEN_309; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _GEN_311 = 3'h7 == exReg_predOp_1_s2Addr[2:0] ? predReg_7 : _GEN_310; // @[Execute.scala 215:62 Execute.scala 215:62]
  wire  _T_308 = _GEN_311 ^ exReg_predOp_1_s2Addr[3]; // @[Execute.scala 215:62]
  wire  _T_309 = _T_305 | _T_308; // @[Execute.scala 74:22]
  wire  _T_310 = _T_305 & _T_308; // @[Execute.scala 75:23]
  wire  _T_311 = _T_305 ^ _T_308; // @[Execute.scala 76:23]
  wire  _T_313 = ~_T_309; // @[Execute.scala 77:19]
  wire  _T_315 = 2'h1 == exReg_predOp_1_func ? _T_310 : _T_309; // @[Mux.scala 80:57]
  wire  _T_317 = 2'h2 == exReg_predOp_1_func ? _T_311 : _T_315; // @[Mux.scala 80:57]
  wire  _T_319 = 2'h3 == exReg_predOp_1_func ? _T_313 : _T_317; // @[Mux.scala 80:57]
  wire  _T_322 = exReg_aluOp_1_isCmp ? _T_289 : _T_319; // @[Execute.scala 219:43]
  wire  _GEN_313 = 3'h1 == exReg_predOp_1_dest ? _T_322 : _GEN_255; // @[Execute.scala 219:37 Execute.scala 219:37]
  wire  _GEN_314 = 3'h2 == exReg_predOp_1_dest ? _T_322 : _GEN_256; // @[Execute.scala 219:37 Execute.scala 219:37]
  wire  _GEN_315 = 3'h3 == exReg_predOp_1_dest ? _T_322 : _GEN_257; // @[Execute.scala 219:37 Execute.scala 219:37]
  wire  _GEN_316 = 3'h4 == exReg_predOp_1_dest ? _T_322 : _GEN_258; // @[Execute.scala 219:37 Execute.scala 219:37]
  wire  _GEN_317 = 3'h5 == exReg_predOp_1_dest ? _T_322 : _GEN_259; // @[Execute.scala 219:37 Execute.scala 219:37]
  wire  _GEN_318 = 3'h6 == exReg_predOp_1_dest ? _T_322 : _GEN_260; // @[Execute.scala 219:37 Execute.scala 219:37]
  wire  _GEN_319 = 3'h7 == exReg_predOp_1_dest ? _T_322 : _GEN_261; // @[Execute.scala 219:37 Execute.scala 219:37]
  wire  _GEN_321 = (exReg_aluOp_1_isCmp | exReg_aluOp_1_isPred) & doExecute_1 ? _GEN_313 : _GEN_255; // @[Execute.scala 218:75]
  wire  _GEN_322 = (exReg_aluOp_1_isCmp | exReg_aluOp_1_isPred) & doExecute_1 ? _GEN_314 : _GEN_256; // @[Execute.scala 218:75]
  wire  _GEN_323 = (exReg_aluOp_1_isCmp | exReg_aluOp_1_isPred) & doExecute_1 ? _GEN_315 : _GEN_257; // @[Execute.scala 218:75]
  wire  _GEN_324 = (exReg_aluOp_1_isCmp | exReg_aluOp_1_isPred) & doExecute_1 ? _GEN_316 : _GEN_258; // @[Execute.scala 218:75]
  wire  _GEN_325 = (exReg_aluOp_1_isCmp | exReg_aluOp_1_isPred) & doExecute_1 ? _GEN_317 : _GEN_259; // @[Execute.scala 218:75]
  wire  _GEN_326 = (exReg_aluOp_1_isCmp | exReg_aluOp_1_isPred) & doExecute_1 ? _GEN_318 : _GEN_260; // @[Execute.scala 218:75]
  wire  _GEN_327 = (exReg_aluOp_1_isCmp | exReg_aluOp_1_isPred) & doExecute_1 ? _GEN_319 : _GEN_261; // @[Execute.scala 218:75]
  wire  _T_338 = 4'h8 == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire  _T_339 = 4'h9 == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire  _T_340 = 4'ha == exReg_aluOp_1_func; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_328 = _T_340 ? op_2 : _GEN_268; // @[Conditional.scala 39:67 Execute.scala 257:21]
  wire [31:0] _GEN_329 = _T_339 ? op_2 : _GEN_267; // @[Conditional.scala 39:67 Execute.scala 254:22]
  wire [31:0] _GEN_330 = _T_339 ? _GEN_268 : _GEN_328; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_331 = _T_338 ? op_2 : _GEN_266; // @[Conditional.scala 39:67 Execute.scala 251:21]
  wire [31:0] _GEN_332 = _T_338 ? _GEN_267 : _GEN_329; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_333 = _T_338 ? _GEN_268 : _GEN_330; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_334 = _T_257 ? op_2 : _GEN_265; // @[Conditional.scala 39:67 Execute.scala 248:22]
  wire [31:0] _GEN_335 = _T_257 ? _GEN_266 : _GEN_331; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_336 = _T_257 ? _GEN_267 : _GEN_332; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_337 = _T_257 ? _GEN_268 : _GEN_333; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_338 = _T_250 ? 3'h2 : _GEN_264; // @[Conditional.scala 39:67 Execute.scala 245:22]
  wire [31:0] _GEN_339 = _T_250 ? _GEN_265 : _GEN_334; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_340 = _T_250 ? _GEN_266 : _GEN_335; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_341 = _T_250 ? _GEN_267 : _GEN_336; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_342 = _T_250 ? _GEN_268 : _GEN_337; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_343 = _T_255 ? 3'h1 : _GEN_338; // @[Conditional.scala 39:67 Execute.scala 242:22]
  wire [31:0] _GEN_344 = _T_255 ? _GEN_265 : _GEN_339; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_345 = _T_255 ? _GEN_266 : _GEN_340; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_346 = _T_255 ? _GEN_267 : _GEN_341; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_347 = _T_255 ? _GEN_268 : _GEN_342; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_348 = _T_246 ? op_2 : _GEN_263; // @[Conditional.scala 39:67 Execute.scala 239:20]
  wire [2:0] _GEN_349 = _T_246 ? _GEN_264 : _GEN_343; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_350 = _T_246 ? _GEN_265 : _GEN_344; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_351 = _T_246 ? _GEN_266 : _GEN_345; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_352 = _T_246 ? _GEN_267 : _GEN_346; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_353 = _T_246 ? _GEN_268 : _GEN_347; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_356 = _T_244 ? _GEN_264 : _GEN_349; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_357 = _T_244 ? _GEN_265 : _GEN_350; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_358 = _T_244 ? _GEN_266 : _GEN_351; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_359 = _T_244 ? _GEN_267 : _GEN_352; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_360 = _T_244 ? _GEN_268 : _GEN_353; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_371 = _T_240 ? _GEN_264 : _GEN_356; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_392 = _T_340 ? excOffReg : 32'h0; // @[Conditional.scala 39:67 Execute.scala 289:19 Execute.scala 262:15]
  wire [31:0] _GEN_393 = _T_339 ? excBaseReg : _GEN_392; // @[Conditional.scala 39:67 Execute.scala 286:19]
  wire [31:0] _GEN_394 = _T_338 ? retOffReg : _GEN_393; // @[Conditional.scala 39:67 Execute.scala 283:19]
  wire [31:0] _GEN_395 = _T_257 ? retBaseReg : _GEN_394; // @[Conditional.scala 39:67 Execute.scala 280:19]
  wire [31:0] _GEN_396 = _T_250 ? io_scex_memTop : _GEN_395; // @[Conditional.scala 39:67 Execute.scala 277:19]
  wire [31:0] _GEN_397 = _T_255 ? io_scex_stackTop : _GEN_396; // @[Conditional.scala 39:67 Execute.scala 274:19]
  wire [31:0] _GEN_398 = _T_246 ? mulHiReg : _GEN_397; // @[Conditional.scala 39:67 Execute.scala 271:19]
  wire [31:0] _GEN_399 = _T_244 ? mulLoReg : _GEN_398; // @[Conditional.scala 39:67 Execute.scala 268:19]
  wire [31:0] _GEN_400 = _T_240 ? _T_216 : _GEN_399; // @[Conditional.scala 40:58 Execute.scala 265:19]
  wire [31:0] _T_352 = exReg_aluOp_1_isBCpy ? _T_302 : _GEN_287[31:0]; // @[Execute.scala 297:35]
  wire  _T_358 = exReg_call & doExecute_0; // @[Execute.scala 312:35]
  wire  _T_362 = exReg_xcall & doExecute_0; // @[Execute.scala 316:37]
  wire  _T_366 = exReg_call | exReg_ret | exReg_brcf | exReg_xcall; // @[Execute.scala 322:58]
  wire [31:0] brcfOff = exReg_immOp_0 ? 32'h0 : op_1; // @[Execute.scala 325:20]
  wire  _T_368 = exReg_call | exReg_xcall; // @[Execute.scala 326:36]
  wire [31:0] _T_369 = exReg_xret ? excOffReg : retOffReg; // @[Execute.scala 328:32]
  wire [31:0] _T_370 = exReg_brcf ? brcfOff : _T_369; // @[Execute.scala 327:28]
  wire [31:0] callRetAddr = exReg_call | exReg_xcall ? 32'h0 : _T_370; // @[Execute.scala 326:24]
  wire [31:0] callBase = exReg_immOp_0 ? exReg_callAddr : op_0; // @[Execute.scala 330:21]
  wire [31:0] _T_373 = exReg_xret ? excBaseReg : retBaseReg; // @[Execute.scala 332:28]
  wire [31:0] callRetBase = _T_368 | exReg_brcf ? callBase : _T_373; // @[Execute.scala 331:24]
  wire [31:0] _T_375 = {exReg_base,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_380 = {exReg_relPc,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_433 = {{2'd0}, op_0[31:2]}; // @[Execute.scala 355:50]
  wire [31:0] _T_384 = _GEN_433 - exReg_jmpOp_reloc; // @[Execute.scala 355:50]
  wire [31:0] target = exReg_immOp_0 ? {{2'd0}, exReg_jmpOp_target} : _T_384; // @[Execute.scala 353:19]
  wire [29:0] hi_6 = saveND ? exReg_relPc : io_feex_pc; // @[Execute.scala 382:25]
  wire [31:0] _T_390 = {hi_6,2'h0}; // @[Cat.scala 30:58]
  assign io_brflush = exReg_nonDelayed & exReg_jmpOp_branch & doExecute_0; // @[Execute.scala 357:56]
  assign io_exmem_rd_0_addr = exReg_rdAddr_0; // @[Execute.scala 294:25]
  assign io_exmem_rd_0_data = exReg_aluOp_0_isMFS ? _GEN_277 : _T_226; // @[Execute.scala 296:31]
  assign io_exmem_rd_0_valid = exReg_wrRd_0 & doExecute_0; // @[Execute.scala 295:43]
  assign io_exmem_rd_1_addr = exReg_rdAddr_1; // @[Execute.scala 294:25]
  assign io_exmem_rd_1_data = exReg_aluOp_1_isMFS ? _GEN_400 : _T_352; // @[Execute.scala 296:31]
  assign io_exmem_rd_1_valid = exReg_wrRd_1 & doExecute_1; // @[Execute.scala 295:43]
  assign io_exmem_mem_load = exReg_memOp_load & doExecute_0; // @[Execute.scala 302:41]
  assign io_exmem_mem_store = exReg_memOp_store & doExecute_0; // @[Execute.scala 303:43]
  assign io_exmem_mem_hword = exReg_memOp_hword; // @[Execute.scala 304:22]
  assign io_exmem_mem_byte = exReg_memOp_byte; // @[Execute.scala 305:21]
  assign io_exmem_mem_zext = exReg_memOp_zext; // @[Execute.scala 306:21]
  assign io_exmem_mem_typ = exReg_memOp_typ; // @[Execute.scala 307:20]
  assign io_exmem_mem_addr = op_0 + exReg_immVal_0; // @[Execute.scala 308:30]
  assign io_exmem_mem_data = fwReg_1[0] ? _GEN_120 : _T_44; // @[Execute.scala 125:21]
  assign io_exmem_mem_call = exReg_call & doExecute_0; // @[Execute.scala 312:35]
  assign io_exmem_mem_ret = exReg_ret & doExecute_0; // @[Execute.scala 313:34]
  assign io_exmem_mem_brcf = exReg_brcf & doExecute_0; // @[Execute.scala 314:35]
  assign io_exmem_mem_trap = exReg_trap & doExecute_0; // @[Execute.scala 315:35]
  assign io_exmem_mem_xcall = exReg_xcall & doExecute_0; // @[Execute.scala 316:37]
  assign io_exmem_mem_xret = exReg_xret & doExecute_0; // @[Execute.scala 317:35]
  assign io_exmem_mem_xsrc = exReg_xsrc; // @[Execute.scala 318:21]
  assign io_exmem_mem_illOp = exReg_illOp; // @[Execute.scala 320:22]
  assign io_exmem_mem_nonDelayed = exReg_nonDelayed; // @[Execute.scala 319:27]
  assign io_exmem_base = exReg_base; // @[Execute.scala 361:17]
  assign io_exmem_relPc = exReg_relPc; // @[Execute.scala 362:18]
  assign io_exicache_doCallRet = (_T_366 | exReg_xret) & doExecute_0; // @[Execute.scala 323:47]
  assign io_exicache_callRetBase = {{2'd0}, callRetBase[31:2]}; // @[Execute.scala 366:41]
  assign io_exicache_callRetAddr = {{2'd0}, callRetAddr[31:2]}; // @[Execute.scala 367:41]
  assign io_exfe_doBranch = exReg_jmpOp_branch & doExecute_0; // @[Execute.scala 352:42]
  assign io_exfe_branchPc = target[29:0]; // @[Execute.scala 356:20]
  assign io_exsc_op = exReg_aluOp_1_isMTS & doExecute_1 ? _GEN_371 : _GEN_264; // @[Execute.scala 224:48]
  assign io_exsc_opData = exReg_aluOp_1_isMTS & doExecute_1 ? op_2 : _GEN_253; // @[Execute.scala 224:48 Execute.scala 225:22]
  assign io_exsc_opOff = exReg_immOp_0 ? exReg_immVal_0 : op_0; // @[Execute.scala 195:23]
  always @(posedge clock) begin
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_base <= io_decex_base; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_relPc <= io_decex_relPc;
    end
    if (reset) begin // @[Execute.scala 386:15]
      exReg_pred_0 <= 4'h8; // @[connections.scala 134:10]
    end else if (io_ena) begin // @[Execute.scala 19:16]
      if (io_flush | io_brflush) begin // @[Execute.scala 21:34]
        exReg_pred_0 <= 4'h8; // @[connections.scala 134:10]
      end else begin
        exReg_pred_0 <= io_decex_pred_0; // @[Execute.scala 20:11]
      end
    end
    if (reset) begin // @[Execute.scala 386:15]
      exReg_pred_1 <= 4'h8; // @[connections.scala 134:10]
    end else if (io_ena) begin // @[Execute.scala 19:16]
      if (io_flush | io_brflush) begin // @[Execute.scala 21:34]
        exReg_pred_1 <= 4'h8; // @[connections.scala 134:10]
      end else begin
        exReg_pred_1 <= io_decex_pred_1; // @[Execute.scala 20:11]
      end
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_0_func <= io_decex_aluOp_0_func; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_0_isMul <= io_decex_aluOp_0_isMul; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_0_isCmp <= io_decex_aluOp_0_isCmp; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_0_isPred <= io_decex_aluOp_0_isPred; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_0_isBCpy <= io_decex_aluOp_0_isBCpy; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_0_isMTS <= io_decex_aluOp_0_isMTS; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_0_isMFS <= io_decex_aluOp_0_isMFS; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_1_func <= io_decex_aluOp_1_func; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_1_isCmp <= io_decex_aluOp_1_isCmp; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_1_isPred <= io_decex_aluOp_1_isPred; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_1_isBCpy <= io_decex_aluOp_1_isBCpy; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_1_isMTS <= io_decex_aluOp_1_isMTS; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_aluOp_1_isMFS <= io_decex_aluOp_1_isMFS; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_predOp_0_func <= io_decex_predOp_0_func; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_predOp_0_dest <= io_decex_predOp_0_dest; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_predOp_0_s1Addr <= io_decex_predOp_0_s1Addr; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_predOp_0_s2Addr <= io_decex_predOp_0_s2Addr; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_predOp_1_func <= io_decex_predOp_1_func; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_predOp_1_dest <= io_decex_predOp_1_dest; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_predOp_1_s1Addr <= io_decex_predOp_1_s1Addr; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_predOp_1_s2Addr <= io_decex_predOp_1_s2Addr; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_jmpOp_branch <= io_decex_jmpOp_branch; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_jmpOp_target <= io_decex_jmpOp_target; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_jmpOp_reloc <= io_decex_jmpOp_reloc; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_memOp_load <= io_decex_memOp_load; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_memOp_store <= io_decex_memOp_store; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_memOp_hword <= io_decex_memOp_hword; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_memOp_byte <= io_decex_memOp_byte; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_memOp_zext <= io_decex_memOp_zext; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_memOp_typ <= io_decex_memOp_typ; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_stackOp <= io_decex_stackOp; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_rsData_0 <= io_decex_rsData_0; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_rsData_1 <= io_decex_rsData_1; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_rsData_2 <= io_decex_rsData_2; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_rsData_3 <= io_decex_rsData_3; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_rdAddr_0 <= io_decex_rdAddr_0; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_rdAddr_1 <= io_decex_rdAddr_1; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_immVal_0 <= io_decex_immVal_0; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_immVal_1 <= io_decex_immVal_1; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_immOp_0 <= io_decex_immOp_0; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_wrRd_0 <= io_decex_wrRd_0; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_wrRd_1 <= io_decex_wrRd_1; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_callAddr <= io_decex_callAddr; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_call <= io_decex_call; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_ret <= io_decex_ret; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_brcf <= io_decex_brcf; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_trap <= io_decex_trap; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_xcall <= io_decex_xcall; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_xret <= io_decex_xret; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_xsrc <= io_decex_xsrc; // @[Execute.scala 20:11]
    end
    if (io_ena) begin // @[Execute.scala 19:16]
      exReg_nonDelayed <= io_decex_nonDelayed; // @[Execute.scala 20:11]
    end
    if (reset) begin // @[Execute.scala 386:15]
      exReg_illOp <= 1'h0; // @[connections.scala 135:11]
    end else if (io_ena) begin // @[Execute.scala 19:16]
      if (io_flush | io_brflush) begin // @[Execute.scala 21:34]
        exReg_illOp <= 1'h0; // @[connections.scala 135:11]
      end else begin
        exReg_illOp <= io_decex_illOp; // @[Execute.scala 20:11]
      end
    end
    if (!(~io_ena)) begin // @[Execute.scala 110:18]
      if (io_decex_rsAddr_0 == io_exResult_1_addr & io_exResult_1_valid) begin // @[Execute.scala 98:80]
        fwReg_0 <= 3'h1; // @[Execute.scala 99:18]
      end else if (io_decex_rsAddr_0 == io_exResult_0_addr & io_exResult_0_valid) begin // @[Execute.scala 98:80]
        fwReg_0 <= 3'h1; // @[Execute.scala 99:18]
      end else if (io_decex_rsAddr_0 == io_memResult_1_addr & io_memResult_1_valid) begin // @[Execute.scala 92:82]
        fwReg_0 <= 3'h2; // @[Execute.scala 93:18]
      end else begin
        fwReg_0 <= _GEN_67;
      end
    end
    if (!(~io_ena)) begin // @[Execute.scala 110:18]
      if (io_decex_immOp_0) begin // @[Execute.scala 105:29]
        fwReg_1 <= 3'h4; // @[Execute.scala 106:20]
      end else if (io_decex_rsAddr_1 == io_exResult_1_addr & io_exResult_1_valid) begin // @[Execute.scala 98:80]
        fwReg_1 <= 3'h1; // @[Execute.scala 99:18]
      end else if (io_decex_rsAddr_1 == io_exResult_0_addr & io_exResult_0_valid) begin // @[Execute.scala 98:80]
        fwReg_1 <= 3'h1; // @[Execute.scala 99:18]
      end else begin
        fwReg_1 <= _GEN_77;
      end
    end
    if (!(~io_ena)) begin // @[Execute.scala 110:18]
      if (io_decex_rsAddr_2 == io_exResult_1_addr & io_exResult_1_valid) begin // @[Execute.scala 98:80]
        fwReg_2 <= 3'h1; // @[Execute.scala 99:18]
      end else if (io_decex_rsAddr_2 == io_exResult_0_addr & io_exResult_0_valid) begin // @[Execute.scala 98:80]
        fwReg_2 <= 3'h1; // @[Execute.scala 99:18]
      end else if (io_decex_rsAddr_2 == io_memResult_1_addr & io_memResult_1_valid) begin // @[Execute.scala 92:82]
        fwReg_2 <= 3'h2; // @[Execute.scala 93:18]
      end else begin
        fwReg_2 <= _GEN_83;
      end
    end
    if (!(~io_ena)) begin // @[Execute.scala 110:18]
      if (io_decex_immOp_1) begin // @[Execute.scala 105:29]
        fwReg_3 <= 3'h4; // @[Execute.scala 106:20]
      end else if (io_decex_rsAddr_3 == io_exResult_1_addr & io_exResult_1_valid) begin // @[Execute.scala 98:80]
        fwReg_3 <= 3'h1; // @[Execute.scala 99:18]
      end else if (io_decex_rsAddr_3 == io_exResult_0_addr & io_exResult_0_valid) begin // @[Execute.scala 98:80]
        fwReg_3 <= 3'h1; // @[Execute.scala 99:18]
      end else begin
        fwReg_3 <= _GEN_93;
      end
    end
    if (!(~io_ena)) begin // @[Execute.scala 110:18]
      fwSrcReg_0 <= _GEN_74;
    end
    if (!(~io_ena)) begin // @[Execute.scala 110:18]
      fwSrcReg_1 <= _GEN_82;
    end
    if (!(~io_ena)) begin // @[Execute.scala 110:18]
      fwSrcReg_2 <= _GEN_90;
    end
    if (!(~io_ena)) begin // @[Execute.scala 110:18]
      fwSrcReg_3 <= _GEN_98;
    end
    if (io_ena) begin // @[Execute.scala 114:17]
      memResultDataReg_0 <= io_memResult_0_data; // @[Execute.scala 115:22]
    end
    if (io_ena) begin // @[Execute.scala 114:17]
      memResultDataReg_1 <= io_memResult_1_data; // @[Execute.scala 115:22]
    end
    if (io_ena) begin // @[Execute.scala 114:17]
      exResultDataReg_0 <= io_exResult_0_data; // @[Execute.scala 116:21]
    end
    if (io_ena) begin // @[Execute.scala 114:17]
      exResultDataReg_1 <= io_exResult_1_data; // @[Execute.scala 116:21]
    end
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          predReg_1 <= op_2[1]; // @[Execute.scala 230:24]
        end else begin
          predReg_1 <= _GEN_321;
        end
      end else begin
        predReg_1 <= _GEN_321;
      end
    end
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          predReg_2 <= op_2[2]; // @[Execute.scala 230:24]
        end else begin
          predReg_2 <= _GEN_322;
        end
      end else begin
        predReg_2 <= _GEN_322;
      end
    end
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          predReg_3 <= op_2[3]; // @[Execute.scala 230:24]
        end else begin
          predReg_3 <= _GEN_323;
        end
      end else begin
        predReg_3 <= _GEN_323;
      end
    end
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          predReg_4 <= op_2[4]; // @[Execute.scala 230:24]
        end else begin
          predReg_4 <= _GEN_324;
        end
      end else begin
        predReg_4 <= _GEN_324;
      end
    end
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          predReg_5 <= op_2[5]; // @[Execute.scala 230:24]
        end else begin
          predReg_5 <= _GEN_325;
        end
      end else begin
        predReg_5 <= _GEN_325;
      end
    end
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          predReg_6 <= op_2[6]; // @[Execute.scala 230:24]
        end else begin
          predReg_6 <= _GEN_326;
        end
      end else begin
        predReg_6 <= _GEN_326;
      end
    end
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          predReg_7 <= op_2[7]; // @[Execute.scala 230:24]
        end else begin
          predReg_7 <= _GEN_327;
        end
      end else begin
        predReg_7 <= _GEN_327;
      end
    end
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (_T_358) begin // @[Execute.scala 338:36]
        retBaseReg <= _T_375; // @[Execute.scala 339:16]
      end else if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          retBaseReg <= _GEN_265;
        end else begin
          retBaseReg <= _GEN_357;
        end
      end else begin
        retBaseReg <= _GEN_265;
      end
    end
    if (saveRetOff) begin // @[Execute.scala 381:20]
      retOffReg <= _T_390; // @[Execute.scala 382:15]
    end else if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          retOffReg <= _GEN_266;
        end else begin
          retOffReg <= _GEN_358;
        end
      end else begin
        retOffReg <= _GEN_266;
      end
    end
    saveRetOff <= _T_358 & io_ena; // @[Execute.scala 342:44]
    saveND <= exReg_nonDelayed; // @[Execute.scala 343:10]
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (_T_362) begin // @[Execute.scala 346:37]
        excBaseReg <= _T_375; // @[Execute.scala 347:16]
      end else if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          excBaseReg <= _GEN_267;
        end else begin
          excBaseReg <= _GEN_359;
        end
      end else begin
        excBaseReg <= _GEN_267;
      end
    end
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (_T_362) begin // @[Execute.scala 346:37]
        excOffReg <= _T_380; // @[Execute.scala 348:15]
      end else if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          excOffReg <= _GEN_268;
        end else begin
          excOffReg <= _GEN_360;
        end
      end else begin
        excOffReg <= _GEN_268;
      end
    end
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          mulLoReg <= _GEN_262;
        end else if (_T_244) begin // @[Conditional.scala 39:67]
          mulLoReg <= op_2; // @[Execute.scala 236:20]
        end else begin
          mulLoReg <= _GEN_262;
        end
      end else begin
        mulLoReg <= _GEN_262;
      end
    end
    if (!(_T_35)) begin // @[Execute.scala 370:17]
      if (exReg_aluOp_1_isMTS & doExecute_1) begin // @[Execute.scala 224:48]
        if (_T_240) begin // @[Conditional.scala 40:58]
          mulHiReg <= _GEN_263;
        end else if (_T_244) begin // @[Conditional.scala 39:67]
          mulHiReg <= _GEN_263;
        end else begin
          mulHiReg <= _GEN_348;
        end
      end else begin
        mulHiReg <= _GEN_263;
      end
    end
    if (io_ena) begin // @[Execute.scala 165:16]
      mulLLReg <= _T_74; // @[Execute.scala 177:14]
    end
    if (io_ena) begin // @[Execute.scala 165:16]
      mulLHReg <= _T_78; // @[Execute.scala 178:14]
    end
    if (io_ena) begin // @[Execute.scala 165:16]
      mulHLReg <= _T_82; // @[Execute.scala 179:14]
    end
    mulHHReg <= _GEN_151[31:0];
    if (io_ena) begin // @[Execute.scala 165:16]
      mulPipeReg <= exReg_aluOp_0_isMul & doExecute_0; // @[Execute.scala 166:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  exReg_base = _RAND_0[29:0];
  _RAND_1 = {1{`RANDOM}};
  exReg_relPc = _RAND_1[29:0];
  _RAND_2 = {1{`RANDOM}};
  exReg_pred_0 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  exReg_pred_1 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  exReg_aluOp_0_func = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  exReg_aluOp_0_isMul = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  exReg_aluOp_0_isCmp = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  exReg_aluOp_0_isPred = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  exReg_aluOp_0_isBCpy = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  exReg_aluOp_0_isMTS = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  exReg_aluOp_0_isMFS = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  exReg_aluOp_1_func = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  exReg_aluOp_1_isCmp = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  exReg_aluOp_1_isPred = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  exReg_aluOp_1_isBCpy = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  exReg_aluOp_1_isMTS = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  exReg_aluOp_1_isMFS = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  exReg_predOp_0_func = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  exReg_predOp_0_dest = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  exReg_predOp_0_s1Addr = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  exReg_predOp_0_s2Addr = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  exReg_predOp_1_func = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  exReg_predOp_1_dest = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  exReg_predOp_1_s1Addr = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  exReg_predOp_1_s2Addr = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  exReg_jmpOp_branch = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  exReg_jmpOp_target = _RAND_26[29:0];
  _RAND_27 = {1{`RANDOM}};
  exReg_jmpOp_reloc = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  exReg_memOp_load = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  exReg_memOp_store = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  exReg_memOp_hword = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  exReg_memOp_byte = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  exReg_memOp_zext = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  exReg_memOp_typ = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  exReg_stackOp = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  exReg_rsData_0 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  exReg_rsData_1 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  exReg_rsData_2 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  exReg_rsData_3 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  exReg_rdAddr_0 = _RAND_39[4:0];
  _RAND_40 = {1{`RANDOM}};
  exReg_rdAddr_1 = _RAND_40[4:0];
  _RAND_41 = {1{`RANDOM}};
  exReg_immVal_0 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  exReg_immVal_1 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  exReg_immOp_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  exReg_wrRd_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  exReg_wrRd_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  exReg_callAddr = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  exReg_call = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  exReg_ret = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  exReg_brcf = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  exReg_trap = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  exReg_xcall = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  exReg_xret = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  exReg_xsrc = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  exReg_nonDelayed = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  exReg_illOp = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  fwReg_0 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  fwReg_1 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  fwReg_2 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  fwReg_3 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  fwSrcReg_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  fwSrcReg_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  fwSrcReg_2 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  fwSrcReg_3 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  memResultDataReg_0 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  memResultDataReg_1 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  exResultDataReg_0 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  exResultDataReg_1 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  predReg_1 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  predReg_2 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  predReg_3 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  predReg_4 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  predReg_5 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  predReg_6 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  predReg_7 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  retBaseReg = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  retOffReg = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  saveRetOff = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  saveND = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  excBaseReg = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  excOffReg = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  mulLoReg = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  mulHiReg = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  mulLLReg = _RAND_83[31:0];
  _RAND_84 = {2{`RANDOM}};
  mulLHReg = _RAND_84[32:0];
  _RAND_85 = {2{`RANDOM}};
  mulHLReg = _RAND_85[32:0];
  _RAND_86 = {1{`RANDOM}};
  mulHHReg = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  mulPipeReg = _RAND_87[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Memory(
  input         clock,
  input         reset,
  output        io_ena_out,
  input         io_ena_in,
  output        io_flush,
  input  [4:0]  io_exmem_rd_0_addr,
  input  [31:0] io_exmem_rd_0_data,
  input         io_exmem_rd_0_valid,
  input  [4:0]  io_exmem_rd_1_addr,
  input  [31:0] io_exmem_rd_1_data,
  input         io_exmem_rd_1_valid,
  input         io_exmem_mem_load,
  input         io_exmem_mem_store,
  input         io_exmem_mem_hword,
  input         io_exmem_mem_byte,
  input         io_exmem_mem_zext,
  input  [1:0]  io_exmem_mem_typ,
  input  [31:0] io_exmem_mem_addr,
  input  [31:0] io_exmem_mem_data,
  input         io_exmem_mem_call,
  input         io_exmem_mem_ret,
  input         io_exmem_mem_brcf,
  input         io_exmem_mem_trap,
  input         io_exmem_mem_xcall,
  input         io_exmem_mem_xret,
  input  [4:0]  io_exmem_mem_xsrc,
  input         io_exmem_mem_illOp,
  input         io_exmem_mem_nonDelayed,
  input  [29:0] io_exmem_base,
  input  [29:0] io_exmem_relPc,
  output [4:0]  io_memwb_rd_0_addr,
  output [31:0] io_memwb_rd_0_data,
  output        io_memwb_rd_0_valid,
  output [4:0]  io_memwb_rd_1_addr,
  output [31:0] io_memwb_rd_1_data,
  output        io_memwb_rd_1_valid,
  output        io_memfe_doCallRet,
  output        io_memfe_store,
  output [31:0] io_memfe_addr,
  output [31:0] io_memfe_data,
  output [4:0]  io_exResult_0_addr,
  output [31:0] io_exResult_0_data,
  output        io_exResult_0_valid,
  output [4:0]  io_exResult_1_addr,
  output [31:0] io_exResult_1_data,
  output        io_exResult_1_valid,
  output [2:0]  io_localInOut_M_Cmd,
  output [31:0] io_localInOut_M_Addr,
  output [31:0] io_localInOut_M_Data,
  output [3:0]  io_localInOut_M_ByteEn,
  input  [1:0]  io_localInOut_S_Resp,
  input  [31:0] io_localInOut_S_Data,
  output [2:0]  io_globalInOut_M_Cmd,
  output [31:0] io_globalInOut_M_Addr,
  output [31:0] io_globalInOut_M_Data,
  output [3:0]  io_globalInOut_M_ByteEn,
  output [1:0]  io_globalInOut_M_AddrSpace,
  input  [1:0]  io_globalInOut_S_Resp,
  input  [31:0] io_globalInOut_S_Data,
  input         io_icacheIllMem,
  input         io_scacheIllMem,
  output        io_exc_call,
  output        io_exc_ret,
  output [4:0]  io_exc_src,
  output        io_exc_exc,
  output [29:0] io_exc_excBase,
  output [29:0] io_exc_excAddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] memReg_rd_0_addr; // @[Memory.scala 21:19]
  reg [31:0] memReg_rd_0_data; // @[Memory.scala 21:19]
  reg  memReg_rd_0_valid; // @[Memory.scala 21:19]
  reg [4:0] memReg_rd_1_addr; // @[Memory.scala 21:19]
  reg [31:0] memReg_rd_1_data; // @[Memory.scala 21:19]
  reg  memReg_rd_1_valid; // @[Memory.scala 21:19]
  reg  memReg_mem_load; // @[Memory.scala 21:19]
  reg  memReg_mem_hword; // @[Memory.scala 21:19]
  reg  memReg_mem_byte; // @[Memory.scala 21:19]
  reg  memReg_mem_zext; // @[Memory.scala 21:19]
  reg [1:0] memReg_mem_typ; // @[Memory.scala 21:19]
  reg [31:0] memReg_mem_addr; // @[Memory.scala 21:19]
  reg  memReg_mem_call; // @[Memory.scala 21:19]
  reg  memReg_mem_ret; // @[Memory.scala 21:19]
  reg  memReg_mem_brcf; // @[Memory.scala 21:19]
  reg  memReg_mem_trap; // @[Memory.scala 21:19]
  reg  memReg_mem_xcall; // @[Memory.scala 21:19]
  reg  memReg_mem_xret; // @[Memory.scala 21:19]
  reg [4:0] memReg_mem_xsrc; // @[Memory.scala 21:19]
  reg  memReg_mem_illOp; // @[Memory.scala 21:19]
  reg  memReg_mem_nonDelayed; // @[Memory.scala 21:19]
  reg [29:0] memReg_base; // @[Memory.scala 21:19]
  reg [29:0] memReg_relPc; // @[Memory.scala 21:19]
  wire  _T_1 = io_globalInOut_S_Resp == 2'h3; // @[Memory.scala 25:39]
  wire  _T_2 = io_localInOut_S_Resp == 2'h3 | _T_1; // @[Memory.scala 24:54]
  wire  _T_3 = _T_2 | io_icacheIllMem; // @[Memory.scala 25:55]
  wire  illMem = _T_3 | io_scacheIllMem; // @[Memory.scala 26:33]
  reg  illMemReg; // @[Memory.scala 27:22]
  wire  _T_6 = memReg_mem_call | memReg_mem_ret | memReg_mem_brcf; // @[Memory.scala 31:52]
  wire  _T_8 = (_T_6 | memReg_mem_xret) & memReg_mem_nonDelayed; // @[Memory.scala 32:54]
  wire  _T_9 = memReg_mem_xcall | memReg_mem_trap | _T_8; // @[Memory.scala 30:52]
  wire  _T_10 = _T_9 | memReg_mem_illOp; // @[Memory.scala 32:80]
  wire  flush = _T_10 | illMemReg; // @[Memory.scala 33:33]
  reg  mayStallReg; // @[Memory.scala 37:28]
  wire  _T_11 = io_localInOut_S_Resp == 2'h1; // @[Memory.scala 38:38]
  wire  _T_13 = _T_11 | io_globalInOut_S_Resp == 2'h1; // @[Memory.scala 39:17]
  wire  enable = _T_13 | ~mayStallReg; // @[Memory.scala 40:17]
  wire  _T_15 = enable & io_ena_in; // @[Memory.scala 44:15]
  wire  _GEN_11 = flush ? 1'h0 : io_exmem_mem_load | io_exmem_mem_store; // @[Memory.scala 47:17 Memory.scala 49:19 Memory.scala 46:17]
  wire  _GEN_40 = enable & io_ena_in ? _GEN_11 : mayStallReg; // @[Memory.scala 44:29 Memory.scala 37:28]
  wire  _GEN_41 = illMem ? 1'h0 : _GEN_40; // @[Memory.scala 52:16 Memory.scala 53:19]
  wire [7:0] _GEN_49 = io_exmem_mem_addr[1] ? io_exmem_mem_data[7:0] : io_exmem_mem_data[7:0]; // @[Memory.scala 92:52 Memory.scala 93:17 Memory.scala 82:15]
  wire [7:0] _GEN_50 = io_exmem_mem_addr[1] ? io_exmem_mem_data[15:8] : io_exmem_mem_data[15:8]; // @[Memory.scala 92:52 Memory.scala 94:17 Memory.scala 82:15]
  wire [3:0] _GEN_51 = io_exmem_mem_addr[1] ? 4'h3 : 4'hf; // @[Memory.scala 92:52 Memory.scala 95:14 Memory.scala 85:10]
  wire [7:0] _GEN_52 = ~io_exmem_mem_addr[1] ? io_exmem_mem_data[7:0] : io_exmem_mem_data[23:16]; // @[Memory.scala 88:47 Memory.scala 89:17 Memory.scala 82:15]
  wire [7:0] _GEN_53 = ~io_exmem_mem_addr[1] ? io_exmem_mem_data[15:8] : io_exmem_mem_data[31:24]; // @[Memory.scala 88:47 Memory.scala 90:17 Memory.scala 82:15]
  wire [3:0] _GEN_54 = ~io_exmem_mem_addr[1] ? 4'hc : _GEN_51; // @[Memory.scala 88:47 Memory.scala 91:14]
  wire [7:0] _GEN_55 = ~io_exmem_mem_addr[1] ? io_exmem_mem_data[7:0] : _GEN_49; // @[Memory.scala 88:47 Memory.scala 82:15]
  wire [7:0] _GEN_56 = ~io_exmem_mem_addr[1] ? io_exmem_mem_data[15:8] : _GEN_50; // @[Memory.scala 88:47 Memory.scala 82:15]
  wire [7:0] _GEN_57 = io_exmem_mem_hword ? _GEN_52 : io_exmem_mem_data[23:16]; // @[Memory.scala 87:28 Memory.scala 82:15]
  wire [7:0] _GEN_58 = io_exmem_mem_hword ? _GEN_53 : io_exmem_mem_data[31:24]; // @[Memory.scala 87:28 Memory.scala 82:15]
  wire [3:0] _GEN_59 = io_exmem_mem_hword ? _GEN_54 : 4'hf; // @[Memory.scala 87:28 Memory.scala 85:10]
  wire [7:0] _GEN_60 = io_exmem_mem_hword ? _GEN_55 : io_exmem_mem_data[7:0]; // @[Memory.scala 87:28 Memory.scala 82:15]
  wire [7:0] _GEN_61 = io_exmem_mem_hword ? _GEN_56 : io_exmem_mem_data[15:8]; // @[Memory.scala 87:28 Memory.scala 82:15]
  wire  _T_36 = 2'h0 == io_exmem_mem_addr[1:0]; // @[Conditional.scala 37:30]
  wire  _T_38 = 2'h1 == io_exmem_mem_addr[1:0]; // @[Conditional.scala 37:30]
  wire  _T_40 = 2'h2 == io_exmem_mem_addr[1:0]; // @[Conditional.scala 37:30]
  wire  _T_42 = 2'h3 == io_exmem_mem_addr[1:0]; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_62 = _T_42 ? io_exmem_mem_data[7:0] : _GEN_60; // @[Conditional.scala 39:67 Memory.scala 114:19]
  wire [3:0] _GEN_63 = _T_42 ? 4'h1 : _GEN_59; // @[Conditional.scala 39:67 Memory.scala 115:16]
  wire [7:0] _GEN_64 = _T_40 ? io_exmem_mem_data[7:0] : _GEN_61; // @[Conditional.scala 39:67 Memory.scala 110:19]
  wire [3:0] _GEN_65 = _T_40 ? 4'h2 : _GEN_63; // @[Conditional.scala 39:67 Memory.scala 111:16]
  wire [7:0] _GEN_66 = _T_40 ? _GEN_60 : _GEN_62; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_67 = _T_38 ? io_exmem_mem_data[7:0] : _GEN_57; // @[Conditional.scala 39:67 Memory.scala 106:19]
  wire [3:0] _GEN_68 = _T_38 ? 4'h4 : _GEN_65; // @[Conditional.scala 39:67 Memory.scala 107:16]
  wire [7:0] _GEN_69 = _T_38 ? _GEN_61 : _GEN_64; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_70 = _T_38 ? _GEN_60 : _GEN_66; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_71 = _T_36 ? io_exmem_mem_data[7:0] : _GEN_58; // @[Conditional.scala 40:58 Memory.scala 102:19]
  wire [3:0] _GEN_72 = _T_36 ? 4'h8 : _GEN_68; // @[Conditional.scala 40:58 Memory.scala 103:16]
  wire [7:0] _GEN_73 = _T_36 ? _GEN_57 : _GEN_67; // @[Conditional.scala 40:58]
  wire [7:0] _GEN_74 = _T_36 ? _GEN_61 : _GEN_69; // @[Conditional.scala 40:58]
  wire [7:0] _GEN_75 = _T_36 ? _GEN_60 : _GEN_70; // @[Conditional.scala 40:58]
  wire [7:0] wrData_3 = io_exmem_mem_byte ? _GEN_71 : _GEN_58; // @[Memory.scala 99:27]
  wire [7:0] wrData_2 = io_exmem_mem_byte ? _GEN_73 : _GEN_57; // @[Memory.scala 99:27]
  wire [7:0] wrData_1 = io_exmem_mem_byte ? _GEN_74 : _GEN_61; // @[Memory.scala 99:27]
  wire [7:0] wrData_0 = io_exmem_mem_byte ? _GEN_75 : _GEN_60; // @[Memory.scala 99:27]
  wire [2:0] _T_48 = {1'h0,io_exmem_mem_load,io_exmem_mem_store}; // @[Memory.scala 123:49]
  wire [2:0] cmd = _T_15 & ~flush ? _T_48 : 3'h0; // @[Memory.scala 122:16]
  wire [29:0] hi = io_exmem_mem_addr[31:2]; // @[Memory.scala 127:48]
  wire [15:0] lo = {wrData_1,wrData_0}; // @[Cat.scala 30:58]
  wire [15:0] hi_1 = {wrData_3,wrData_2}; // @[Cat.scala 30:58]
  wire [1:0] _T_59 = io_exmem_mem_typ == 2'h2 ? 2'h2 : 2'h3; // @[Memory.scala 136:40]
  wire [31:0] _T_63 = memReg_mem_typ == 2'h1 ? io_localInOut_S_Data : io_globalInOut_S_Data; // @[Memory.scala 150:33]
  wire [7:0] rdData_0 = _T_63[7:0]; // @[Memory.scala 142:24]
  wire [7:0] rdData_1 = _T_63[15:8]; // @[Memory.scala 142:24]
  wire [7:0] rdData_2 = _T_63[23:16]; // @[Memory.scala 142:24]
  wire [7:0] rdData_3 = _T_63[31:24]; // @[Memory.scala 142:24]
  wire [15:0] lo_2 = {rdData_1,rdData_0}; // @[Cat.scala 30:58]
  wire [15:0] hi_4 = {rdData_3,rdData_2}; // @[Cat.scala 30:58]
  wire [31:0] _T_69 = {rdData_3,rdData_2,rdData_1,rdData_0}; // @[Cat.scala 30:58]
  wire [7:0] _T_72 = 2'h1 == memReg_mem_addr[1:0] ? rdData_2 : rdData_3; // @[Mux.scala 80:57]
  wire [7:0] _T_74 = 2'h2 == memReg_mem_addr[1:0] ? rdData_1 : _T_72; // @[Mux.scala 80:57]
  wire [7:0] bval = 2'h3 == memReg_mem_addr[1:0] ? rdData_0 : _T_74; // @[Mux.scala 80:57]
  wire [15:0] hval = ~memReg_mem_addr[1] ? hi_4 : lo_2; // @[Memory.scala 164:17]
  wire [23:0] _T_82 = bval[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  wire [23:0] _T_83 = memReg_mem_zext ? 24'h0 : _T_82; // @[Memory.scala 170:16]
  wire [31:0] _T_84 = {_T_83,bval}; // @[Memory.scala 172:66]
  wire [31:0] _GEN_81 = memReg_mem_byte ? _T_84 : _T_69; // @[Memory.scala 169:25 Memory.scala 170:10 Memory.scala 155:8]
  wire [15:0] _T_87 = hval[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_88 = memReg_mem_zext ? 16'h0 : _T_87; // @[Memory.scala 175:16]
  wire [31:0] _T_89 = {_T_88,hval}; // @[Memory.scala 177:70]
  wire [31:0] dout = memReg_mem_hword ? _T_89 : _GEN_81; // @[Memory.scala 174:26 Memory.scala 175:10]
  wire  _T_93 = _T_6 | memReg_mem_xcall; // @[Memory.scala 186:79]
  wire [4:0] _T_101 = illMemReg ? 5'h1 : memReg_mem_xsrc; // @[Memory.scala 206:24]
  wire [29:0] _T_104 = memReg_relPc + 30'h1; // @[Memory.scala 209:55]
  assign io_ena_out = _T_13 | ~mayStallReg; // @[Memory.scala 40:17]
  assign io_flush = _T_10 | illMemReg; // @[Memory.scala 33:33]
  assign io_memwb_rd_0_addr = memReg_rd_0_addr; // @[Memory.scala 181:15]
  assign io_memwb_rd_0_data = memReg_mem_load ? dout : memReg_rd_0_data; // @[Memory.scala 183:29]
  assign io_memwb_rd_0_valid = memReg_rd_0_valid; // @[Memory.scala 181:15]
  assign io_memwb_rd_1_addr = memReg_rd_1_addr; // @[Memory.scala 181:15]
  assign io_memwb_rd_1_data = memReg_rd_1_data; // @[Memory.scala 181:15]
  assign io_memwb_rd_1_valid = memReg_rd_1_valid; // @[Memory.scala 181:15]
  assign io_memfe_doCallRet = _T_93 | memReg_mem_xret; // @[Memory.scala 187:43]
  assign io_memfe_store = io_localInOut_M_Cmd == 3'h1; // @[Memory.scala 192:41]
  assign io_memfe_addr = io_exmem_mem_addr; // @[Memory.scala 193:17]
  assign io_memfe_data = {hi_1,lo}; // @[Cat.scala 30:58]
  assign io_exResult_0_addr = io_exmem_rd_0_addr; // @[Memory.scala 197:15]
  assign io_exResult_0_data = io_exmem_rd_0_data; // @[Memory.scala 197:15]
  assign io_exResult_0_valid = io_exmem_rd_0_valid; // @[Memory.scala 197:15]
  assign io_exResult_1_addr = io_exmem_rd_1_addr; // @[Memory.scala 197:15]
  assign io_exResult_1_data = io_exmem_rd_1_data; // @[Memory.scala 197:15]
  assign io_exResult_1_valid = io_exmem_rd_1_valid; // @[Memory.scala 197:15]
  assign io_localInOut_M_Cmd = io_exmem_mem_typ == 2'h1 ? cmd : 3'h0; // @[Memory.scala 126:29]
  assign io_localInOut_M_Addr = {hi,2'h0}; // @[Cat.scala 30:58]
  assign io_localInOut_M_Data = {hi_1,lo}; // @[Cat.scala 30:58]
  assign io_localInOut_M_ByteEn = io_exmem_mem_byte ? _GEN_72 : _GEN_59; // @[Memory.scala 99:27]
  assign io_globalInOut_M_Cmd = io_exmem_mem_typ != 2'h1 ? cmd : 3'h0; // @[Memory.scala 131:30]
  assign io_globalInOut_M_Addr = {hi,2'h0}; // @[Cat.scala 30:58]
  assign io_globalInOut_M_Data = {hi_1,lo}; // @[Cat.scala 30:58]
  assign io_globalInOut_M_ByteEn = io_exmem_mem_byte ? _GEN_72 : _GEN_59; // @[Memory.scala 99:27]
  assign io_globalInOut_M_AddrSpace = io_exmem_mem_typ == 2'h0 ? 2'h0 : _T_59; // @[Memory.scala 135:36]
  assign io_exc_call = memReg_mem_xcall; // @[Memory.scala 200:15]
  assign io_exc_ret = memReg_mem_xret; // @[Memory.scala 201:14]
  assign io_exc_src = memReg_mem_illOp ? 5'h0 : _T_101; // @[Memory.scala 205:20]
  assign io_exc_exc = memReg_mem_trap | memReg_mem_illOp | illMemReg; // @[Memory.scala 203:53]
  assign io_exc_excBase = memReg_base; // @[Memory.scala 208:18]
  assign io_exc_excAddr = memReg_mem_trap ? _T_104 : memReg_relPc; // @[Memory.scala 209:24]
  always @(posedge clock) begin
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_rd_0_addr <= io_exmem_rd_0_addr; // @[Memory.scala 45:12]
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_rd_0_data <= io_exmem_rd_0_data; // @[Memory.scala 45:12]
    end
    if (reset) begin // @[Memory.scala 215:15]
      memReg_rd_0_valid <= 1'h0; // @[connections.scala 172:11]
    end else if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      if (flush) begin // @[Memory.scala 47:17]
        memReg_rd_0_valid <= 1'h0; // @[connections.scala 172:11]
      end else begin
        memReg_rd_0_valid <= io_exmem_rd_0_valid; // @[Memory.scala 45:12]
      end
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_rd_1_addr <= io_exmem_rd_1_addr; // @[Memory.scala 45:12]
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_rd_1_data <= io_exmem_rd_1_data; // @[Memory.scala 45:12]
    end
    if (reset) begin // @[Memory.scala 215:15]
      memReg_rd_1_valid <= 1'h0; // @[connections.scala 172:11]
    end else if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      if (flush) begin // @[Memory.scala 47:17]
        memReg_rd_1_valid <= 1'h0; // @[connections.scala 172:11]
      end else begin
        memReg_rd_1_valid <= io_exmem_rd_1_valid; // @[Memory.scala 45:12]
      end
    end
    if (reset) begin // @[Memory.scala 215:15]
      memReg_mem_load <= 1'h0; // @[connections.scala 198:10]
    end else if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      if (flush) begin // @[Memory.scala 47:17]
        memReg_mem_load <= 1'h0; // @[connections.scala 198:10]
      end else begin
        memReg_mem_load <= io_exmem_mem_load; // @[Memory.scala 45:12]
      end
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_mem_hword <= io_exmem_mem_hword; // @[Memory.scala 45:12]
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_mem_byte <= io_exmem_mem_byte; // @[Memory.scala 45:12]
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_mem_zext <= io_exmem_mem_zext; // @[Memory.scala 45:12]
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_mem_typ <= io_exmem_mem_typ; // @[Memory.scala 45:12]
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_mem_addr <= io_exmem_mem_addr; // @[Memory.scala 45:12]
    end
    if (reset) begin // @[Memory.scala 215:15]
      memReg_mem_call <= 1'h0; // @[connections.scala 200:10]
    end else if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      if (flush) begin // @[Memory.scala 47:17]
        memReg_mem_call <= 1'h0; // @[connections.scala 200:10]
      end else begin
        memReg_mem_call <= io_exmem_mem_call; // @[Memory.scala 45:12]
      end
    end
    if (reset) begin // @[Memory.scala 215:15]
      memReg_mem_ret <= 1'h0; // @[connections.scala 201:9]
    end else if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      if (flush) begin // @[Memory.scala 47:17]
        memReg_mem_ret <= 1'h0; // @[connections.scala 201:9]
      end else begin
        memReg_mem_ret <= io_exmem_mem_ret; // @[Memory.scala 45:12]
      end
    end
    if (reset) begin // @[Memory.scala 215:15]
      memReg_mem_brcf <= 1'h0; // @[connections.scala 202:10]
    end else if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      if (flush) begin // @[Memory.scala 47:17]
        memReg_mem_brcf <= 1'h0; // @[connections.scala 202:10]
      end else begin
        memReg_mem_brcf <= io_exmem_mem_brcf; // @[Memory.scala 45:12]
      end
    end
    if (reset) begin // @[Memory.scala 215:15]
      memReg_mem_trap <= 1'h0; // @[connections.scala 203:10]
    end else if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      if (flush) begin // @[Memory.scala 47:17]
        memReg_mem_trap <= 1'h0; // @[connections.scala 203:10]
      end else begin
        memReg_mem_trap <= io_exmem_mem_trap; // @[Memory.scala 45:12]
      end
    end
    if (reset) begin // @[Memory.scala 215:15]
      memReg_mem_xcall <= 1'h0; // @[connections.scala 204:11]
    end else if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      if (flush) begin // @[Memory.scala 47:17]
        memReg_mem_xcall <= 1'h0; // @[connections.scala 204:11]
      end else begin
        memReg_mem_xcall <= io_exmem_mem_xcall; // @[Memory.scala 45:12]
      end
    end
    if (reset) begin // @[Memory.scala 215:15]
      memReg_mem_xret <= 1'h0; // @[connections.scala 205:10]
    end else if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      if (flush) begin // @[Memory.scala 47:17]
        memReg_mem_xret <= 1'h0; // @[connections.scala 205:10]
      end else begin
        memReg_mem_xret <= io_exmem_mem_xret; // @[Memory.scala 45:12]
      end
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_mem_xsrc <= io_exmem_mem_xsrc; // @[Memory.scala 45:12]
    end
    if (reset) begin // @[Memory.scala 215:15]
      memReg_mem_illOp <= 1'h0; // @[connections.scala 206:11]
    end else if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      if (flush) begin // @[Memory.scala 47:17]
        memReg_mem_illOp <= 1'h0; // @[connections.scala 206:11]
      end else begin
        memReg_mem_illOp <= io_exmem_mem_illOp; // @[Memory.scala 45:12]
      end
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_mem_nonDelayed <= io_exmem_mem_nonDelayed; // @[Memory.scala 45:12]
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_base <= io_exmem_base; // @[Memory.scala 45:12]
    end
    if (enable & io_ena_in) begin // @[Memory.scala 44:29]
      memReg_relPc <= io_exmem_relPc; // @[Memory.scala 45:12]
    end
    illMemReg <= _T_3 | io_scacheIllMem; // @[Memory.scala 26:33]
    if (reset) begin // @[Memory.scala 37:28]
      mayStallReg <= 1'h0; // @[Memory.scala 37:28]
    end else if (~io_ena_in) begin // @[Memory.scala 60:21]
      if (io_localInOut_S_Resp != 2'h0 | io_globalInOut_S_Resp != 2'h0) begin // @[Memory.scala 61:92]
        mayStallReg <= 1'h0; // @[Memory.scala 62:19]
      end else begin
        mayStallReg <= _GEN_41;
      end
    end else begin
      mayStallReg <= _GEN_41;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_rd_0_addr = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  memReg_rd_0_data = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_rd_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  memReg_rd_1_addr = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_rd_1_data = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  memReg_rd_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  memReg_mem_load = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  memReg_mem_hword = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  memReg_mem_byte = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  memReg_mem_zext = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  memReg_mem_typ = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  memReg_mem_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  memReg_mem_call = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  memReg_mem_ret = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  memReg_mem_brcf = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  memReg_mem_trap = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  memReg_mem_xcall = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  memReg_mem_xret = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  memReg_mem_xsrc = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  memReg_mem_illOp = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  memReg_mem_nonDelayed = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  memReg_base = _RAND_21[29:0];
  _RAND_22 = {1{`RANDOM}};
  memReg_relPc = _RAND_22[29:0];
  _RAND_23 = {1{`RANDOM}};
  illMemReg = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  mayStallReg = _RAND_24[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WriteBack(
  input  [4:0]  io_memwb_rd_0_addr,
  input  [31:0] io_memwb_rd_0_data,
  input         io_memwb_rd_0_valid,
  input  [4:0]  io_memwb_rd_1_addr,
  input  [31:0] io_memwb_rd_1_data,
  input         io_memwb_rd_1_valid,
  output [4:0]  io_rfWrite_0_addr,
  output [31:0] io_rfWrite_0_data,
  output        io_rfWrite_0_valid,
  output [4:0]  io_rfWrite_1_addr,
  output [31:0] io_rfWrite_1_data,
  output        io_rfWrite_1_valid,
  output [4:0]  io_memResult_0_addr,
  output [31:0] io_memResult_0_data,
  output        io_memResult_0_valid,
  output [4:0]  io_memResult_1_addr,
  output [31:0] io_memResult_1_data,
  output        io_memResult_1_valid
);
  assign io_rfWrite_0_addr = io_memwb_rd_0_addr; // @[WriteBack.scala 21:14]
  assign io_rfWrite_0_data = io_memwb_rd_0_data; // @[WriteBack.scala 21:14]
  assign io_rfWrite_0_valid = io_memwb_rd_0_valid; // @[WriteBack.scala 21:14]
  assign io_rfWrite_1_addr = io_memwb_rd_1_addr; // @[WriteBack.scala 21:14]
  assign io_rfWrite_1_data = io_memwb_rd_1_data; // @[WriteBack.scala 21:14]
  assign io_rfWrite_1_valid = io_memwb_rd_1_valid; // @[WriteBack.scala 21:14]
  assign io_memResult_0_addr = io_memwb_rd_0_addr; // @[WriteBack.scala 23:16]
  assign io_memResult_0_data = io_memwb_rd_0_data; // @[WriteBack.scala 23:16]
  assign io_memResult_0_valid = io_memwb_rd_0_valid; // @[WriteBack.scala 23:16]
  assign io_memResult_1_addr = io_memwb_rd_1_addr; // @[WriteBack.scala 23:16]
  assign io_memResult_1_data = io_memwb_rd_1_data; // @[WriteBack.scala 23:16]
  assign io_memResult_1_valid = io_memwb_rd_1_valid; // @[WriteBack.scala 23:16]
endmodule
module Exceptions(
  input         clock,
  input         reset,
  input         io_ena,
  input  [2:0]  io_ocp_M_Cmd,
  input  [31:0] io_ocp_M_Addr,
  input  [31:0] io_ocp_M_Data,
  output [1:0]  io_ocp_S_Resp,
  output [31:0] io_ocp_S_Data,
  input         io_intrs_0,
  input         io_intrs_1,
  input         io_intrs_2,
  input         io_intrs_3,
  input         io_intrs_4,
  input         io_intrs_5,
  output        io_excdec_exc,
  output [29:0] io_excdec_excBase,
  output [29:0] io_excdec_excAddr,
  output        io_excdec_intr,
  output [31:0] io_excdec_addr,
  output [4:0]  io_excdec_src,
  output        io_excdec_local,
  input         io_memexc_call,
  input         io_memexc_ret,
  input  [4:0]  io_memexc_src,
  input         io_memexc_exc,
  input  [29:0] io_memexc_excBase,
  input  [29:0] io_memexc_excAddr,
  output        io_invalICache,
  output        io_invalDCache
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] vec [0:31];
  wire [31:0] vec_MPORT_data;
  wire [4:0] vec_MPORT_addr;
  wire [31:0] vec_MPORT_1_data;
  wire [4:0] vec_MPORT_1_addr;
  wire  vec_MPORT_1_mask;
  wire  vec_MPORT_1_en;
  reg [31:0] vecDup [0:31];
  wire [31:0] vecDup_MPORT_3_data;
  wire [4:0] vecDup_MPORT_3_addr;
  wire [31:0] vecDup_MPORT_2_data;
  wire [4:0] vecDup_MPORT_2_addr;
  wire  vecDup_MPORT_2_mask;
  wire  vecDup_MPORT_2_en;
  reg [2:0] masterReg_Cmd; // @[Exceptions.scala 21:26]
  reg [31:0] masterReg_Addr; // @[Exceptions.scala 21:26]
  reg [31:0] masterReg_Data; // @[Exceptions.scala 21:26]
  reg [31:0] statusReg; // @[Exceptions.scala 23:26]
  reg [31:0] maskReg; // @[Exceptions.scala 24:22]
  reg [31:0] sourceReg; // @[Exceptions.scala 25:22]
  wire  intrEna = statusReg[0]; // @[Exceptions.scala 27:26]
  wire  superMode = statusReg[1]; // @[Exceptions.scala 28:28]
  reg  localModeReg; // @[Exceptions.scala 30:29]
  reg  sleepReg; // @[Exceptions.scala 39:25]
  reg  excPendReg_0; // @[Exceptions.scala 43:28]
  reg  excPendReg_1; // @[Exceptions.scala 43:28]
  reg  excPendReg_2; // @[Exceptions.scala 43:28]
  reg  excPendReg_3; // @[Exceptions.scala 43:28]
  reg  excPendReg_4; // @[Exceptions.scala 43:28]
  reg  excPendReg_5; // @[Exceptions.scala 43:28]
  reg  excPendReg_6; // @[Exceptions.scala 43:28]
  reg  excPendReg_7; // @[Exceptions.scala 43:28]
  reg  excPendReg_8; // @[Exceptions.scala 43:28]
  reg  excPendReg_9; // @[Exceptions.scala 43:28]
  reg  excPendReg_10; // @[Exceptions.scala 43:28]
  reg  excPendReg_11; // @[Exceptions.scala 43:28]
  reg  excPendReg_12; // @[Exceptions.scala 43:28]
  reg  excPendReg_13; // @[Exceptions.scala 43:28]
  reg  excPendReg_14; // @[Exceptions.scala 43:28]
  reg  excPendReg_15; // @[Exceptions.scala 43:28]
  reg  excPendReg_16; // @[Exceptions.scala 43:28]
  reg  excPendReg_17; // @[Exceptions.scala 43:28]
  reg  excPendReg_18; // @[Exceptions.scala 43:28]
  reg  excPendReg_19; // @[Exceptions.scala 43:28]
  reg  excPendReg_20; // @[Exceptions.scala 43:28]
  reg  excPendReg_21; // @[Exceptions.scala 43:28]
  reg  excPendReg_22; // @[Exceptions.scala 43:28]
  reg  excPendReg_23; // @[Exceptions.scala 43:28]
  reg  excPendReg_24; // @[Exceptions.scala 43:28]
  reg  excPendReg_25; // @[Exceptions.scala 43:28]
  reg  excPendReg_26; // @[Exceptions.scala 43:28]
  reg  excPendReg_27; // @[Exceptions.scala 43:28]
  reg  excPendReg_28; // @[Exceptions.scala 43:28]
  reg  excPendReg_29; // @[Exceptions.scala 43:28]
  reg  excPendReg_30; // @[Exceptions.scala 43:28]
  reg  excPendReg_31; // @[Exceptions.scala 43:28]
  reg  intrPendReg_16; // @[Exceptions.scala 45:28]
  reg  intrPendReg_17; // @[Exceptions.scala 45:28]
  reg  intrPendReg_18; // @[Exceptions.scala 45:28]
  reg  intrPendReg_19; // @[Exceptions.scala 45:28]
  reg  intrPendReg_20; // @[Exceptions.scala 45:28]
  reg  intrPendReg_21; // @[Exceptions.scala 45:28]
  wire  _T_2 = masterReg_Cmd == 3'h2; // @[Exceptions.scala 61:22]
  wire  _T_4 = 6'h0 == masterReg_Addr[7:2]; // @[Conditional.scala 37:30]
  wire  _T_5 = 6'h1 == masterReg_Addr[7:2]; // @[Conditional.scala 37:30]
  wire  _T_6 = 6'h3 == masterReg_Addr[7:2]; // @[Conditional.scala 37:30]
  wire  _T_7 = 6'h2 == masterReg_Addr[7:2]; // @[Conditional.scala 37:30]
  wire [31:0] _T_8 = {8'h0,2'h0,intrPendReg_21,intrPendReg_20,intrPendReg_19,intrPendReg_18,intrPendReg_17,
    intrPendReg_16,16'h0}; // @[Exceptions.scala 68:58]
  wire  _T_9 = 6'h5 == masterReg_Addr[7:2]; // @[Conditional.scala 37:30]
  wire [31:0] _T_10 = {localModeReg,31'h0}; // @[Exceptions.scala 69:59]
  wire [31:0] _GEN_0 = _T_9 ? _T_10 : 32'h0; // @[Conditional.scala 39:67 Exceptions.scala 69:43 Exceptions.scala 51:17]
  wire [31:0] _GEN_1 = _T_7 ? _T_8 : _GEN_0; // @[Conditional.scala 39:67 Exceptions.scala 68:43]
  wire [31:0] _GEN_2 = _T_6 ? sourceReg : _GEN_1; // @[Conditional.scala 39:67 Exceptions.scala 67:43]
  wire [31:0] _GEN_3 = _T_5 ? maskReg : _GEN_2; // @[Conditional.scala 39:67 Exceptions.scala 66:43]
  wire [31:0] _GEN_4 = _T_4 ? statusReg : _GEN_3; // @[Conditional.scala 40:58 Exceptions.scala 65:43]
  wire [31:0] _GEN_8 = masterReg_Addr[7] ? vec_MPORT_data : _GEN_4; // @[Exceptions.scala 71:59 Exceptions.scala 72:21]
  wire [1:0] _GEN_9 = masterReg_Cmd == 3'h2 ? 2'h1 : 2'h0; // @[Exceptions.scala 61:37 Exceptions.scala 62:19 Exceptions.scala 50:17]
  wire  _T_14 = masterReg_Cmd == 3'h1; // @[Exceptions.scala 77:22]
  wire [31:0] _GEN_14 = superMode ? masterReg_Data : statusReg; // @[Exceptions.scala 33:22 Exceptions.scala 80:48 Exceptions.scala 23:26]
  wire [1:0] _GEN_15 = superMode ? 2'h1 : 2'h3; // @[Exceptions.scala 33:22 Exceptions.scala 78:19 Exceptions.scala 33:58]
  wire [31:0] _GEN_17 = superMode ? masterReg_Data : sourceReg; // @[Exceptions.scala 33:22 Exceptions.scala 82:48 Exceptions.scala 25:22]
  wire  _GEN_34 = superMode ? intrPendReg_16 & masterReg_Data[16] : intrPendReg_16; // @[Exceptions.scala 33:22 Exceptions.scala 86:25 Exceptions.scala 47:12]
  wire  _GEN_35 = superMode ? intrPendReg_17 & masterReg_Data[17] : intrPendReg_17; // @[Exceptions.scala 33:22 Exceptions.scala 86:25 Exceptions.scala 47:12]
  wire  _GEN_36 = superMode ? intrPendReg_18 & masterReg_Data[18] : intrPendReg_18; // @[Exceptions.scala 33:22 Exceptions.scala 86:25 Exceptions.scala 47:12]
  wire  _GEN_37 = superMode ? intrPendReg_19 & masterReg_Data[19] : intrPendReg_19; // @[Exceptions.scala 33:22 Exceptions.scala 86:25 Exceptions.scala 47:12]
  wire  _GEN_38 = superMode ? intrPendReg_20 & masterReg_Data[20] : intrPendReg_20; // @[Exceptions.scala 33:22 Exceptions.scala 86:25 Exceptions.scala 47:12]
  wire  _GEN_39 = superMode ? intrPendReg_21 & masterReg_Data[21] : intrPendReg_21; // @[Exceptions.scala 33:22 Exceptions.scala 86:25 Exceptions.scala 47:12]
  wire  _T_84 = 6'h4 == masterReg_Addr[7:2]; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_50 = superMode ? 2'h0 : 2'h3; // @[Exceptions.scala 33:22 Exceptions.scala 92:25 Exceptions.scala 33:58]
  wire  _GEN_51 = superMode | sleepReg; // @[Exceptions.scala 33:22 Exceptions.scala 93:20 Exceptions.scala 39:25]
  wire  _GEN_52 = superMode & masterReg_Data[0]; // @[Exceptions.scala 33:22 Exceptions.scala 98:26 Exceptions.scala 58:18]
  wire  _GEN_53 = superMode & masterReg_Data[1]; // @[Exceptions.scala 33:22 Exceptions.scala 99:26 Exceptions.scala 57:18]
  wire  _GEN_54 = superMode ? localModeReg ^ masterReg_Data[31] : localModeReg; // @[Exceptions.scala 33:22 Exceptions.scala 100:24 Exceptions.scala 30:29]
  wire  _GEN_57 = _T_9 ? _GEN_54 : localModeReg; // @[Conditional.scala 39:67 Exceptions.scala 30:29]
  wire [1:0] _GEN_58 = _T_9 ? _GEN_15 : 2'h1; // @[Conditional.scala 39:67 Exceptions.scala 78:19]
  wire [1:0] _GEN_59 = _T_84 ? _GEN_50 : _GEN_58; // @[Conditional.scala 39:67]
  wire  _GEN_60 = _T_84 ? _GEN_51 : sleepReg; // @[Conditional.scala 39:67 Exceptions.scala 39:25]
  wire  _GEN_61 = _T_84 ? 1'h0 : _T_9 & _GEN_52; // @[Conditional.scala 39:67 Exceptions.scala 58:18]
  wire  _GEN_62 = _T_84 ? 1'h0 : _T_9 & _GEN_53; // @[Conditional.scala 39:67 Exceptions.scala 57:18]
  wire  _GEN_63 = _T_84 ? localModeReg : _GEN_57; // @[Conditional.scala 39:67 Exceptions.scala 30:29]
  wire  _GEN_80 = _T_7 ? _GEN_34 : intrPendReg_16; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_81 = _T_7 ? _GEN_35 : intrPendReg_17; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_82 = _T_7 ? _GEN_36 : intrPendReg_18; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_83 = _T_7 ? _GEN_37 : intrPendReg_19; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_84 = _T_7 ? _GEN_38 : intrPendReg_20; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_85 = _T_7 ? _GEN_39 : intrPendReg_21; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire [1:0] _GEN_96 = _T_7 ? _GEN_15 : _GEN_59; // @[Conditional.scala 39:67]
  wire  _GEN_97 = _T_7 ? sleepReg : _GEN_60; // @[Conditional.scala 39:67 Exceptions.scala 39:25]
  wire  _GEN_98 = _T_7 ? 1'h0 : _GEN_61; // @[Conditional.scala 39:67 Exceptions.scala 58:18]
  wire  _GEN_99 = _T_7 ? 1'h0 : _GEN_62; // @[Conditional.scala 39:67 Exceptions.scala 57:18]
  wire  _GEN_100 = _T_7 ? localModeReg : _GEN_63; // @[Conditional.scala 39:67 Exceptions.scala 30:29]
  wire [31:0] _GEN_101 = _T_6 ? _GEN_17 : sourceReg; // @[Conditional.scala 39:67 Exceptions.scala 25:22]
  wire [1:0] _GEN_102 = _T_6 ? _GEN_15 : _GEN_96; // @[Conditional.scala 39:67]
  wire  _GEN_119 = _T_6 ? intrPendReg_16 : _GEN_80; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_120 = _T_6 ? intrPendReg_17 : _GEN_81; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_121 = _T_6 ? intrPendReg_18 : _GEN_82; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_122 = _T_6 ? intrPendReg_19 : _GEN_83; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_123 = _T_6 ? intrPendReg_20 : _GEN_84; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_124 = _T_6 ? intrPendReg_21 : _GEN_85; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_135 = _T_6 ? sleepReg : _GEN_97; // @[Conditional.scala 39:67 Exceptions.scala 39:25]
  wire  _GEN_136 = _T_6 ? 1'h0 : _GEN_98; // @[Conditional.scala 39:67 Exceptions.scala 58:18]
  wire  _GEN_137 = _T_6 ? 1'h0 : _GEN_99; // @[Conditional.scala 39:67 Exceptions.scala 57:18]
  wire  _GEN_138 = _T_6 ? localModeReg : _GEN_100; // @[Conditional.scala 39:67 Exceptions.scala 30:29]
  wire [1:0] _GEN_140 = _T_5 ? _GEN_15 : _GEN_102; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_141 = _T_5 ? sourceReg : _GEN_101; // @[Conditional.scala 39:67 Exceptions.scala 25:22]
  wire  _GEN_158 = _T_5 ? intrPendReg_16 : _GEN_119; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_159 = _T_5 ? intrPendReg_17 : _GEN_120; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_160 = _T_5 ? intrPendReg_18 : _GEN_121; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_161 = _T_5 ? intrPendReg_19 : _GEN_122; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_162 = _T_5 ? intrPendReg_20 : _GEN_123; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_163 = _T_5 ? intrPendReg_21 : _GEN_124; // @[Conditional.scala 39:67 Exceptions.scala 47:12]
  wire  _GEN_174 = _T_5 ? sleepReg : _GEN_135; // @[Conditional.scala 39:67 Exceptions.scala 39:25]
  wire  _GEN_175 = _T_5 ? 1'h0 : _GEN_136; // @[Conditional.scala 39:67 Exceptions.scala 58:18]
  wire  _GEN_176 = _T_5 ? 1'h0 : _GEN_137; // @[Conditional.scala 39:67 Exceptions.scala 57:18]
  wire [31:0] _GEN_178 = _T_4 ? _GEN_14 : statusReg; // @[Conditional.scala 40:58 Exceptions.scala 23:26]
  wire [1:0] _GEN_179 = _T_4 ? _GEN_15 : _GEN_140; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_181 = _T_4 ? sourceReg : _GEN_141; // @[Conditional.scala 40:58 Exceptions.scala 25:22]
  wire  _GEN_198 = _T_4 ? intrPendReg_16 : _GEN_158; // @[Conditional.scala 40:58 Exceptions.scala 47:12]
  wire  _GEN_199 = _T_4 ? intrPendReg_17 : _GEN_159; // @[Conditional.scala 40:58 Exceptions.scala 47:12]
  wire  _GEN_200 = _T_4 ? intrPendReg_18 : _GEN_160; // @[Conditional.scala 40:58 Exceptions.scala 47:12]
  wire  _GEN_201 = _T_4 ? intrPendReg_19 : _GEN_161; // @[Conditional.scala 40:58 Exceptions.scala 47:12]
  wire  _GEN_202 = _T_4 ? intrPendReg_20 : _GEN_162; // @[Conditional.scala 40:58 Exceptions.scala 47:12]
  wire  _GEN_203 = _T_4 ? intrPendReg_21 : _GEN_163; // @[Conditional.scala 40:58 Exceptions.scala 47:12]
  wire  _GEN_215 = _T_4 ? 1'h0 : _GEN_175; // @[Conditional.scala 40:58 Exceptions.scala 58:18]
  wire  _GEN_216 = _T_4 ? 1'h0 : _GEN_176; // @[Conditional.scala 40:58 Exceptions.scala 57:18]
  wire [1:0] _GEN_224 = superMode ? _GEN_179 : 2'h3; // @[Exceptions.scala 33:22 Exceptions.scala 33:58]
  wire  _GEN_227 = masterReg_Addr[7] & superMode; // @[Exceptions.scala 104:59]
  wire [1:0] _GEN_231 = masterReg_Addr[7] ? _GEN_224 : _GEN_179; // @[Exceptions.scala 104:59]
  wire [1:0] _GEN_232 = masterReg_Cmd == 3'h1 ? _GEN_231 : _GEN_9; // @[Exceptions.scala 77:37]
  wire [31:0] _GEN_233 = masterReg_Cmd == 3'h1 ? _GEN_178 : statusReg; // @[Exceptions.scala 77:37 Exceptions.scala 23:26]
  wire [31:0] _GEN_235 = masterReg_Cmd == 3'h1 ? _GEN_181 : sourceReg; // @[Exceptions.scala 77:37 Exceptions.scala 25:22]
  wire  _GEN_252 = masterReg_Cmd == 3'h1 ? _GEN_198 : intrPendReg_16; // @[Exceptions.scala 77:37 Exceptions.scala 47:12]
  wire  _GEN_253 = masterReg_Cmd == 3'h1 ? _GEN_199 : intrPendReg_17; // @[Exceptions.scala 77:37 Exceptions.scala 47:12]
  wire  _GEN_254 = masterReg_Cmd == 3'h1 ? _GEN_200 : intrPendReg_18; // @[Exceptions.scala 77:37 Exceptions.scala 47:12]
  wire  _GEN_255 = masterReg_Cmd == 3'h1 ? _GEN_201 : intrPendReg_19; // @[Exceptions.scala 77:37 Exceptions.scala 47:12]
  wire  _GEN_256 = masterReg_Cmd == 3'h1 ? _GEN_202 : intrPendReg_20; // @[Exceptions.scala 77:37 Exceptions.scala 47:12]
  wire  _GEN_257 = masterReg_Cmd == 3'h1 ? _GEN_203 : intrPendReg_21; // @[Exceptions.scala 77:37 Exceptions.scala 47:12]
  wire  _GEN_278 = 5'h0 == io_memexc_src ? 1'h0 : excPendReg_0; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_279 = 5'h1 == io_memexc_src ? 1'h0 : excPendReg_1; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_280 = 5'h2 == io_memexc_src ? 1'h0 : excPendReg_2; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_281 = 5'h3 == io_memexc_src ? 1'h0 : excPendReg_3; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_282 = 5'h4 == io_memexc_src ? 1'h0 : excPendReg_4; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_283 = 5'h5 == io_memexc_src ? 1'h0 : excPendReg_5; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_284 = 5'h6 == io_memexc_src ? 1'h0 : excPendReg_6; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_285 = 5'h7 == io_memexc_src ? 1'h0 : excPendReg_7; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_286 = 5'h8 == io_memexc_src ? 1'h0 : excPendReg_8; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_287 = 5'h9 == io_memexc_src ? 1'h0 : excPendReg_9; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_288 = 5'ha == io_memexc_src ? 1'h0 : excPendReg_10; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_289 = 5'hb == io_memexc_src ? 1'h0 : excPendReg_11; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_290 = 5'hc == io_memexc_src ? 1'h0 : excPendReg_12; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_291 = 5'hd == io_memexc_src ? 1'h0 : excPendReg_13; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_292 = 5'he == io_memexc_src ? 1'h0 : excPendReg_14; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_293 = 5'hf == io_memexc_src ? 1'h0 : excPendReg_15; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_294 = 5'h10 == io_memexc_src ? 1'h0 : excPendReg_16; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_295 = 5'h11 == io_memexc_src ? 1'h0 : excPendReg_17; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_296 = 5'h12 == io_memexc_src ? 1'h0 : excPendReg_18; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_297 = 5'h13 == io_memexc_src ? 1'h0 : excPendReg_19; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_298 = 5'h14 == io_memexc_src ? 1'h0 : excPendReg_20; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_299 = 5'h15 == io_memexc_src ? 1'h0 : excPendReg_21; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_300 = 5'h16 == io_memexc_src ? 1'h0 : excPendReg_22; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_301 = 5'h17 == io_memexc_src ? 1'h0 : excPendReg_23; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_302 = 5'h18 == io_memexc_src ? 1'h0 : excPendReg_24; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_303 = 5'h19 == io_memexc_src ? 1'h0 : excPendReg_25; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_304 = 5'h1a == io_memexc_src ? 1'h0 : excPendReg_26; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_305 = 5'h1b == io_memexc_src ? 1'h0 : excPendReg_27; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_306 = 5'h1c == io_memexc_src ? 1'h0 : excPendReg_28; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_307 = 5'h1d == io_memexc_src ? 1'h0 : excPendReg_29; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_308 = 5'h1e == io_memexc_src ? 1'h0 : excPendReg_30; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_309 = 5'h1f == io_memexc_src ? 1'h0 : excPendReg_31; // @[Exceptions.scala 114:28 Exceptions.scala 114:28 Exceptions.scala 46:11]
  wire  _GEN_326 = 5'h10 == io_memexc_src ? 1'h0 : _GEN_252; // @[Exceptions.scala 115:29 Exceptions.scala 115:29]
  wire  _GEN_327 = 5'h11 == io_memexc_src ? 1'h0 : _GEN_253; // @[Exceptions.scala 115:29 Exceptions.scala 115:29]
  wire  _GEN_328 = 5'h12 == io_memexc_src ? 1'h0 : _GEN_254; // @[Exceptions.scala 115:29 Exceptions.scala 115:29]
  wire  _GEN_329 = 5'h13 == io_memexc_src ? 1'h0 : _GEN_255; // @[Exceptions.scala 115:29 Exceptions.scala 115:29]
  wire  _GEN_330 = 5'h14 == io_memexc_src ? 1'h0 : _GEN_256; // @[Exceptions.scala 115:29 Exceptions.scala 115:29]
  wire  _GEN_331 = 5'h15 == io_memexc_src ? 1'h0 : _GEN_257; // @[Exceptions.scala 115:29 Exceptions.scala 115:29]
  wire [33:0] _GEN_560 = {statusReg, 2'h0}; // @[Exceptions.scala 119:31]
  wire [34:0] _T_94 = {{1'd0}, _GEN_560}; // @[Exceptions.scala 119:31]
  wire [34:0] _T_95 = _T_94 | 35'h2; // @[Exceptions.scala 119:43]
  wire [34:0] _GEN_343 = io_ena ? _T_95 : {{3'd0}, _GEN_233}; // @[Exceptions.scala 116:18 Exceptions.scala 119:17]
  wire  _GEN_344 = io_memexc_call ? _GEN_278 : excPendReg_0; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_345 = io_memexc_call ? _GEN_279 : excPendReg_1; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_346 = io_memexc_call ? _GEN_280 : excPendReg_2; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_347 = io_memexc_call ? _GEN_281 : excPendReg_3; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_348 = io_memexc_call ? _GEN_282 : excPendReg_4; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_349 = io_memexc_call ? _GEN_283 : excPendReg_5; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_350 = io_memexc_call ? _GEN_284 : excPendReg_6; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_351 = io_memexc_call ? _GEN_285 : excPendReg_7; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_352 = io_memexc_call ? _GEN_286 : excPendReg_8; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_353 = io_memexc_call ? _GEN_287 : excPendReg_9; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_354 = io_memexc_call ? _GEN_288 : excPendReg_10; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_355 = io_memexc_call ? _GEN_289 : excPendReg_11; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_356 = io_memexc_call ? _GEN_290 : excPendReg_12; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_357 = io_memexc_call ? _GEN_291 : excPendReg_13; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_358 = io_memexc_call ? _GEN_292 : excPendReg_14; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_359 = io_memexc_call ? _GEN_293 : excPendReg_15; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_360 = io_memexc_call ? _GEN_294 : excPendReg_16; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_361 = io_memexc_call ? _GEN_295 : excPendReg_17; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_362 = io_memexc_call ? _GEN_296 : excPendReg_18; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_363 = io_memexc_call ? _GEN_297 : excPendReg_19; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_364 = io_memexc_call ? _GEN_298 : excPendReg_20; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_365 = io_memexc_call ? _GEN_299 : excPendReg_21; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_366 = io_memexc_call ? _GEN_300 : excPendReg_22; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_367 = io_memexc_call ? _GEN_301 : excPendReg_23; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_368 = io_memexc_call ? _GEN_302 : excPendReg_24; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_369 = io_memexc_call ? _GEN_303 : excPendReg_25; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_370 = io_memexc_call ? _GEN_304 : excPendReg_26; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_371 = io_memexc_call ? _GEN_305 : excPendReg_27; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_372 = io_memexc_call ? _GEN_306 : excPendReg_28; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_373 = io_memexc_call ? _GEN_307 : excPendReg_29; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_374 = io_memexc_call ? _GEN_308 : excPendReg_30; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_375 = io_memexc_call ? _GEN_309 : excPendReg_31; // @[Exceptions.scala 113:24 Exceptions.scala 46:11]
  wire  _GEN_392 = io_memexc_call ? _GEN_326 : _GEN_252; // @[Exceptions.scala 113:24]
  wire  _GEN_393 = io_memexc_call ? _GEN_327 : _GEN_253; // @[Exceptions.scala 113:24]
  wire  _GEN_394 = io_memexc_call ? _GEN_328 : _GEN_254; // @[Exceptions.scala 113:24]
  wire  _GEN_395 = io_memexc_call ? _GEN_329 : _GEN_255; // @[Exceptions.scala 113:24]
  wire  _GEN_396 = io_memexc_call ? _GEN_330 : _GEN_256; // @[Exceptions.scala 113:24]
  wire  _GEN_397 = io_memexc_call ? _GEN_331 : _GEN_257; // @[Exceptions.scala 113:24]
  wire [34:0] _GEN_409 = io_memexc_call ? _GEN_343 : {{3'd0}, _GEN_233}; // @[Exceptions.scala 113:24]
  wire [31:0] _T_96 = {{2'd0}, statusReg[31:2]}; // @[Exceptions.scala 126:30]
  wire [34:0] _GEN_410 = io_ena ? {{3'd0}, _T_96} : _GEN_409; // @[Exceptions.scala 124:18 Exceptions.scala 126:17]
  wire [34:0] _GEN_411 = io_memexc_ret ? _GEN_410 : _GEN_409; // @[Exceptions.scala 123:23]
  reg  REG; // @[Exceptions.scala 132:17]
  wire  intrPend_16 = REG | _GEN_392; // @[Exceptions.scala 132:32 Exceptions.scala 133:22]
  reg  REG_1; // @[Exceptions.scala 132:17]
  wire  intrPend_17 = REG_1 | _GEN_393; // @[Exceptions.scala 132:32 Exceptions.scala 133:22]
  reg  REG_2; // @[Exceptions.scala 132:17]
  wire  intrPend_18 = REG_2 | _GEN_394; // @[Exceptions.scala 132:32 Exceptions.scala 133:22]
  reg  REG_3; // @[Exceptions.scala 132:17]
  wire  intrPend_19 = REG_3 | _GEN_395; // @[Exceptions.scala 132:32 Exceptions.scala 133:22]
  reg  REG_4; // @[Exceptions.scala 132:17]
  wire  intrPend_20 = REG_4 | _GEN_396; // @[Exceptions.scala 132:32 Exceptions.scala 133:22]
  reg  REG_5; // @[Exceptions.scala 132:17]
  wire  intrPend_21 = REG_5 | _GEN_397; // @[Exceptions.scala 132:32 Exceptions.scala 133:22]
  reg [29:0] excBaseReg; // @[Exceptions.scala 138:23]
  reg [29:0] excAddrReg; // @[Exceptions.scala 139:23]
  wire  _GEN_428 = 5'h0 == io_memexc_src | _GEN_344; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_429 = 5'h1 == io_memexc_src | _GEN_345; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_430 = 5'h2 == io_memexc_src | _GEN_346; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_431 = 5'h3 == io_memexc_src | _GEN_347; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_432 = 5'h4 == io_memexc_src | _GEN_348; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_433 = 5'h5 == io_memexc_src | _GEN_349; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_434 = 5'h6 == io_memexc_src | _GEN_350; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_435 = 5'h7 == io_memexc_src | _GEN_351; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_436 = 5'h8 == io_memexc_src | _GEN_352; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_437 = 5'h9 == io_memexc_src | _GEN_353; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_438 = 5'ha == io_memexc_src | _GEN_354; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_439 = 5'hb == io_memexc_src | _GEN_355; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_440 = 5'hc == io_memexc_src | _GEN_356; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_441 = 5'hd == io_memexc_src | _GEN_357; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_442 = 5'he == io_memexc_src | _GEN_358; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_443 = 5'hf == io_memexc_src | _GEN_359; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_444 = 5'h10 == io_memexc_src | _GEN_360; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_445 = 5'h11 == io_memexc_src | _GEN_361; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_446 = 5'h12 == io_memexc_src | _GEN_362; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_447 = 5'h13 == io_memexc_src | _GEN_363; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_448 = 5'h14 == io_memexc_src | _GEN_364; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_449 = 5'h15 == io_memexc_src | _GEN_365; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_450 = 5'h16 == io_memexc_src | _GEN_366; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_451 = 5'h17 == io_memexc_src | _GEN_367; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_452 = 5'h18 == io_memexc_src | _GEN_368; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_453 = 5'h19 == io_memexc_src | _GEN_369; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_454 = 5'h1a == io_memexc_src | _GEN_370; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_455 = 5'h1b == io_memexc_src | _GEN_371; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_456 = 5'h1c == io_memexc_src | _GEN_372; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_457 = 5'h1d == io_memexc_src | _GEN_373; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_458 = 5'h1e == io_memexc_src | _GEN_374; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  _GEN_459 = 5'h1f == io_memexc_src | _GEN_375; // @[Exceptions.scala 141:28 Exceptions.scala 141:28]
  wire  excPend_0 = io_memexc_exc ? _GEN_428 : _GEN_344; // @[Exceptions.scala 140:23]
  wire  excPend_1 = io_memexc_exc ? _GEN_429 : _GEN_345; // @[Exceptions.scala 140:23]
  wire  excPend_2 = io_memexc_exc ? _GEN_430 : _GEN_346; // @[Exceptions.scala 140:23]
  wire  excPend_3 = io_memexc_exc ? _GEN_431 : _GEN_347; // @[Exceptions.scala 140:23]
  wire  excPend_4 = io_memexc_exc ? _GEN_432 : _GEN_348; // @[Exceptions.scala 140:23]
  wire  excPend_5 = io_memexc_exc ? _GEN_433 : _GEN_349; // @[Exceptions.scala 140:23]
  wire  excPend_6 = io_memexc_exc ? _GEN_434 : _GEN_350; // @[Exceptions.scala 140:23]
  wire  excPend_7 = io_memexc_exc ? _GEN_435 : _GEN_351; // @[Exceptions.scala 140:23]
  wire  excPend_8 = io_memexc_exc ? _GEN_436 : _GEN_352; // @[Exceptions.scala 140:23]
  wire  excPend_9 = io_memexc_exc ? _GEN_437 : _GEN_353; // @[Exceptions.scala 140:23]
  wire  excPend_10 = io_memexc_exc ? _GEN_438 : _GEN_354; // @[Exceptions.scala 140:23]
  wire  excPend_11 = io_memexc_exc ? _GEN_439 : _GEN_355; // @[Exceptions.scala 140:23]
  wire  excPend_12 = io_memexc_exc ? _GEN_440 : _GEN_356; // @[Exceptions.scala 140:23]
  wire  excPend_13 = io_memexc_exc ? _GEN_441 : _GEN_357; // @[Exceptions.scala 140:23]
  wire  excPend_14 = io_memexc_exc ? _GEN_442 : _GEN_358; // @[Exceptions.scala 140:23]
  wire  excPend_15 = io_memexc_exc ? _GEN_443 : _GEN_359; // @[Exceptions.scala 140:23]
  wire  excPend_16 = io_memexc_exc ? _GEN_444 : _GEN_360; // @[Exceptions.scala 140:23]
  wire  excPend_17 = io_memexc_exc ? _GEN_445 : _GEN_361; // @[Exceptions.scala 140:23]
  wire  excPend_18 = io_memexc_exc ? _GEN_446 : _GEN_362; // @[Exceptions.scala 140:23]
  wire  excPend_19 = io_memexc_exc ? _GEN_447 : _GEN_363; // @[Exceptions.scala 140:23]
  wire  excPend_20 = io_memexc_exc ? _GEN_448 : _GEN_364; // @[Exceptions.scala 140:23]
  wire  excPend_21 = io_memexc_exc ? _GEN_449 : _GEN_365; // @[Exceptions.scala 140:23]
  wire  excPend_22 = io_memexc_exc ? _GEN_450 : _GEN_366; // @[Exceptions.scala 140:23]
  wire  excPend_23 = io_memexc_exc ? _GEN_451 : _GEN_367; // @[Exceptions.scala 140:23]
  wire  excPend_24 = io_memexc_exc ? _GEN_452 : _GEN_368; // @[Exceptions.scala 140:23]
  wire  excPend_25 = io_memexc_exc ? _GEN_453 : _GEN_369; // @[Exceptions.scala 140:23]
  wire  excPend_26 = io_memexc_exc ? _GEN_454 : _GEN_370; // @[Exceptions.scala 140:23]
  wire  excPend_27 = io_memexc_exc ? _GEN_455 : _GEN_371; // @[Exceptions.scala 140:23]
  wire  excPend_28 = io_memexc_exc ? _GEN_456 : _GEN_372; // @[Exceptions.scala 140:23]
  wire  excPend_29 = io_memexc_exc ? _GEN_457 : _GEN_373; // @[Exceptions.scala 140:23]
  wire  excPend_30 = io_memexc_exc ? _GEN_458 : _GEN_374; // @[Exceptions.scala 140:23]
  wire  excPend_31 = io_memexc_exc ? _GEN_459 : _GEN_375; // @[Exceptions.scala 140:23]
  reg [4:0] srcReg; // @[Exceptions.scala 152:23]
  wire [4:0] _GEN_504 = intrPend_21 & maskReg[21] ? 5'h15 : 5'h0; // @[Exceptions.scala 155:51 Exceptions.scala 155:57]
  wire [4:0] _GEN_505 = intrPend_20 & maskReg[20] ? 5'h14 : _GEN_504; // @[Exceptions.scala 155:51 Exceptions.scala 155:57]
  wire [4:0] _GEN_506 = intrPend_19 & maskReg[19] ? 5'h13 : _GEN_505; // @[Exceptions.scala 155:51 Exceptions.scala 155:57]
  wire [4:0] _GEN_507 = intrPend_18 & maskReg[18] ? 5'h12 : _GEN_506; // @[Exceptions.scala 155:51 Exceptions.scala 155:57]
  wire [4:0] _GEN_508 = intrPend_17 & maskReg[17] ? 5'h11 : _GEN_507; // @[Exceptions.scala 155:51 Exceptions.scala 155:57]
  wire [4:0] _GEN_509 = intrPend_16 & maskReg[16] ? 5'h10 : _GEN_508; // @[Exceptions.scala 155:51 Exceptions.scala 155:57]
  wire [4:0] _GEN_526 = excPend_31 ? 5'h1f : _GEN_509; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_527 = excPend_30 ? 5'h1e : _GEN_526; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_528 = excPend_29 ? 5'h1d : _GEN_527; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_529 = excPend_28 ? 5'h1c : _GEN_528; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_530 = excPend_27 ? 5'h1b : _GEN_529; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_531 = excPend_26 ? 5'h1a : _GEN_530; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_532 = excPend_25 ? 5'h19 : _GEN_531; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_533 = excPend_24 ? 5'h18 : _GEN_532; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_534 = excPend_23 ? 5'h17 : _GEN_533; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_535 = excPend_22 ? 5'h16 : _GEN_534; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_536 = excPend_21 ? 5'h15 : _GEN_535; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_537 = excPend_20 ? 5'h14 : _GEN_536; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_538 = excPend_19 ? 5'h13 : _GEN_537; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_539 = excPend_18 ? 5'h12 : _GEN_538; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_540 = excPend_17 ? 5'h11 : _GEN_539; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_541 = excPend_16 ? 5'h10 : _GEN_540; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_542 = excPend_15 ? 5'hf : _GEN_541; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_543 = excPend_14 ? 5'he : _GEN_542; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_544 = excPend_13 ? 5'hd : _GEN_543; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_545 = excPend_12 ? 5'hc : _GEN_544; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_546 = excPend_11 ? 5'hb : _GEN_545; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_547 = excPend_10 ? 5'ha : _GEN_546; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_548 = excPend_9 ? 5'h9 : _GEN_547; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_549 = excPend_8 ? 5'h8 : _GEN_548; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_550 = excPend_7 ? 5'h7 : _GEN_549; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_551 = excPend_6 ? 5'h6 : _GEN_550; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_552 = excPend_5 ? 5'h5 : _GEN_551; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [4:0] _GEN_553 = excPend_4 ? 5'h4 : _GEN_552; // @[Exceptions.scala 158:22 Exceptions.scala 158:28]
  wire [7:0] lo_lo_1 = {excPend_7,excPend_6,excPend_5,excPend_4,excPend_3,excPend_2,excPend_1,excPend_0}; // @[Exceptions.scala 162:29]
  wire [15:0] lo_1 = {excPend_15,excPend_14,excPend_13,excPend_12,excPend_11,excPend_10,excPend_9,excPend_8,lo_lo_1}; // @[Exceptions.scala 162:29]
  wire [7:0] hi_lo_1 = {excPend_23,excPend_22,excPend_21,excPend_20,excPend_19,excPend_18,excPend_17,excPend_16}; // @[Exceptions.scala 162:29]
  wire [31:0] _T_193 = {excPend_31,excPend_30,excPend_29,excPend_28,excPend_27,excPend_26,excPend_25,excPend_24,hi_lo_1,
    lo_1}; // @[Exceptions.scala 162:29]
  reg  exc; // @[Exceptions.scala 162:20]
  wire [31:0] _T_195 = {8'h0,2'h0,intrPend_21,intrPend_20,intrPend_19,intrPend_18,intrPend_17,intrPend_16,16'h0}; // @[Exceptions.scala 163:32]
  wire [31:0] _T_196 = _T_195 & maskReg; // @[Exceptions.scala 163:39]
  reg  intr; // @[Exceptions.scala 163:21]
  wire  _T_198 = intr & intrEna; // @[Exceptions.scala 166:27]
  assign vec_MPORT_addr = masterReg_Addr[6:2];
  assign vec_MPORT_data = vec[vec_MPORT_addr];
  assign vec_MPORT_1_data = masterReg_Data;
  assign vec_MPORT_1_addr = masterReg_Addr[6:2];
  assign vec_MPORT_1_mask = 1'h1;
  assign vec_MPORT_1_en = _T_14 & _GEN_227;
  assign vecDup_MPORT_3_addr = srcReg;
  assign vecDup_MPORT_3_data = vecDup[vecDup_MPORT_3_addr];
  assign vecDup_MPORT_2_data = masterReg_Data;
  assign vecDup_MPORT_2_addr = masterReg_Addr[6:2];
  assign vecDup_MPORT_2_mask = 1'h1;
  assign vecDup_MPORT_2_en = _T_14 & _GEN_227;
  assign io_ocp_S_Resp = sleepReg & (exc | _T_198) ? 2'h1 : _GEN_232; // @[Exceptions.scala 175:61 Exceptions.scala 176:19]
  assign io_ocp_S_Data = masterReg_Cmd == 3'h2 ? _GEN_8 : 32'h0; // @[Exceptions.scala 61:37 Exceptions.scala 51:17]
  assign io_excdec_exc = exc; // @[Exceptions.scala 165:19]
  assign io_excdec_excBase = excBaseReg; // @[Exceptions.scala 171:21]
  assign io_excdec_excAddr = excAddrReg; // @[Exceptions.scala 172:21]
  assign io_excdec_intr = intr & intrEna; // @[Exceptions.scala 166:27]
  assign io_excdec_addr = vecDup_MPORT_3_data; // @[Exceptions.scala 167:19]
  assign io_excdec_src = srcReg; // @[Exceptions.scala 168:19]
  assign io_excdec_local = localModeReg; // @[Exceptions.scala 169:19]
  assign io_invalICache = masterReg_Cmd == 3'h1 & _GEN_216; // @[Exceptions.scala 77:37 Exceptions.scala 57:18]
  assign io_invalDCache = masterReg_Cmd == 3'h1 & _GEN_215; // @[Exceptions.scala 77:37 Exceptions.scala 58:18]
  always @(posedge clock) begin
    if(vec_MPORT_1_en & vec_MPORT_1_mask) begin
      vec[vec_MPORT_1_addr] <= vec_MPORT_1_data;
    end
    if(vecDup_MPORT_2_en & vecDup_MPORT_2_mask) begin
      vecDup[vecDup_MPORT_2_addr] <= vecDup_MPORT_2_data;
    end
    masterReg_Cmd <= io_ocp_M_Cmd; // @[Exceptions.scala 21:26]
    masterReg_Addr <= io_ocp_M_Addr; // @[Exceptions.scala 21:26]
    masterReg_Data <= io_ocp_M_Data; // @[Exceptions.scala 21:26]
    if (reset) begin // @[Exceptions.scala 23:26]
      statusReg <= 32'h2; // @[Exceptions.scala 23:26]
    end else begin
      statusReg <= _GEN_411[31:0];
    end
    if (masterReg_Cmd == 3'h1) begin // @[Exceptions.scala 77:37]
      if (!(_T_4)) begin // @[Conditional.scala 40:58]
        if (_T_5) begin // @[Conditional.scala 39:67]
          if (superMode) begin // @[Exceptions.scala 33:22]
            maskReg <= masterReg_Data; // @[Exceptions.scala 81:46]
          end
        end
      end
    end
    if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (io_ena) begin // @[Exceptions.scala 116:18]
        sourceReg <= {{27'd0}, io_memexc_src}; // @[Exceptions.scala 117:17]
      end else begin
        sourceReg <= _GEN_235;
      end
    end else begin
      sourceReg <= _GEN_235;
    end
    if (reset) begin // @[Exceptions.scala 30:29]
      localModeReg <= 1'h0; // @[Exceptions.scala 30:29]
    end else if (masterReg_Cmd == 3'h1) begin // @[Exceptions.scala 77:37]
      if (!(_T_4)) begin // @[Conditional.scala 40:58]
        if (!(_T_5)) begin // @[Conditional.scala 39:67]
          localModeReg <= _GEN_138;
        end
      end
    end
    if (reset) begin // @[Exceptions.scala 39:25]
      sleepReg <= 1'h0; // @[Exceptions.scala 39:25]
    end else if (sleepReg & (exc | _T_198)) begin // @[Exceptions.scala 175:61]
      sleepReg <= 1'h0; // @[Exceptions.scala 177:14]
    end else if (masterReg_Cmd == 3'h1) begin // @[Exceptions.scala 77:37]
      if (!(_T_4)) begin // @[Conditional.scala 40:58]
        sleepReg <= _GEN_174;
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_0 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_0 <= _GEN_428;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h0 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_0 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_1 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_1 <= _GEN_429;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h1 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_1 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_2 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_2 <= _GEN_430;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h2 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_2 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_3 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_3 <= _GEN_431;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h3 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_3 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_4 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_4 <= _GEN_432;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h4 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_4 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_5 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_5 <= _GEN_433;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h5 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_5 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_6 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_6 <= _GEN_434;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h6 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_6 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_7 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_7 <= _GEN_435;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h7 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_7 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_8 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_8 <= _GEN_436;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h8 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_8 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_9 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_9 <= _GEN_437;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h9 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_9 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_10 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_10 <= _GEN_438;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'ha == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_10 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_11 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_11 <= _GEN_439;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'hb == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_11 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_12 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_12 <= _GEN_440;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'hc == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_12 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_13 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_13 <= _GEN_441;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'hd == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_13 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_14 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_14 <= _GEN_442;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'he == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_14 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_15 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_15 <= _GEN_443;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'hf == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_15 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_16 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_16 <= _GEN_444;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h10 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_16 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_17 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_17 <= _GEN_445;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h11 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_17 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_18 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_18 <= _GEN_446;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h12 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_18 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_19 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_19 <= _GEN_447;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h13 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_19 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_20 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_20 <= _GEN_448;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h14 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_20 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_21 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_21 <= _GEN_449;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h15 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_21 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_22 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_22 <= _GEN_450;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h16 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_22 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_23 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_23 <= _GEN_451;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h17 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_23 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_24 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_24 <= _GEN_452;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h18 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_24 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_25 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_25 <= _GEN_453;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h19 == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_25 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_26 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_26 <= _GEN_454;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h1a == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_26 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_27 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_27 <= _GEN_455;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h1b == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_27 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_28 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_28 <= _GEN_456;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h1c == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_28 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_29 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_29 <= _GEN_457;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h1d == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_29 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_30 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_30 <= _GEN_458;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h1e == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_30 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 43:28]
      excPendReg_31 <= 1'h0; // @[Exceptions.scala 43:28]
    end else if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excPendReg_31 <= _GEN_459;
    end else if (io_memexc_call) begin // @[Exceptions.scala 113:24]
      if (5'h1f == io_memexc_src) begin // @[Exceptions.scala 114:28]
        excPendReg_31 <= 1'h0; // @[Exceptions.scala 114:28]
      end
    end
    if (reset) begin // @[Exceptions.scala 45:28]
      intrPendReg_16 <= 1'h0; // @[Exceptions.scala 45:28]
    end else begin
      intrPendReg_16 <= intrPend_16; // @[Exceptions.scala 148:15]
    end
    if (reset) begin // @[Exceptions.scala 45:28]
      intrPendReg_17 <= 1'h0; // @[Exceptions.scala 45:28]
    end else begin
      intrPendReg_17 <= intrPend_17; // @[Exceptions.scala 148:15]
    end
    if (reset) begin // @[Exceptions.scala 45:28]
      intrPendReg_18 <= 1'h0; // @[Exceptions.scala 45:28]
    end else begin
      intrPendReg_18 <= intrPend_18; // @[Exceptions.scala 148:15]
    end
    if (reset) begin // @[Exceptions.scala 45:28]
      intrPendReg_19 <= 1'h0; // @[Exceptions.scala 45:28]
    end else begin
      intrPendReg_19 <= intrPend_19; // @[Exceptions.scala 148:15]
    end
    if (reset) begin // @[Exceptions.scala 45:28]
      intrPendReg_20 <= 1'h0; // @[Exceptions.scala 45:28]
    end else begin
      intrPendReg_20 <= intrPend_20; // @[Exceptions.scala 148:15]
    end
    if (reset) begin // @[Exceptions.scala 45:28]
      intrPendReg_21 <= 1'h0; // @[Exceptions.scala 45:28]
    end else begin
      intrPendReg_21 <= intrPend_21; // @[Exceptions.scala 148:15]
    end
    REG <= io_intrs_0; // @[Exceptions.scala 132:17]
    REG_1 <= io_intrs_1; // @[Exceptions.scala 132:17]
    REG_2 <= io_intrs_2; // @[Exceptions.scala 132:17]
    REG_3 <= io_intrs_3; // @[Exceptions.scala 132:17]
    REG_4 <= io_intrs_4; // @[Exceptions.scala 132:17]
    REG_5 <= io_intrs_5; // @[Exceptions.scala 132:17]
    if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excBaseReg <= io_memexc_excBase; // @[Exceptions.scala 142:16]
    end
    if (io_memexc_exc) begin // @[Exceptions.scala 140:23]
      excAddrReg <= io_memexc_excAddr; // @[Exceptions.scala 143:16]
    end
    if (excPend_0) begin // @[Exceptions.scala 158:22]
      srcReg <= 5'h0; // @[Exceptions.scala 158:28]
    end else if (excPend_1) begin // @[Exceptions.scala 158:22]
      srcReg <= 5'h1; // @[Exceptions.scala 158:28]
    end else if (excPend_2) begin // @[Exceptions.scala 158:22]
      srcReg <= 5'h2; // @[Exceptions.scala 158:28]
    end else if (excPend_3) begin // @[Exceptions.scala 158:22]
      srcReg <= 5'h3; // @[Exceptions.scala 158:28]
    end else begin
      srcReg <= _GEN_553;
    end
    exc <= _T_193 != 32'h0; // @[Exceptions.scala 162:36]
    intr <= _T_196 != 32'h0; // @[Exceptions.scala 163:50]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    vec[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    vecDup[initvar] = _RAND_1[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  masterReg_Cmd = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  masterReg_Addr = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  masterReg_Data = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  statusReg = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  maskReg = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  sourceReg = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  localModeReg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sleepReg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  excPendReg_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  excPendReg_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  excPendReg_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  excPendReg_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  excPendReg_4 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  excPendReg_5 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  excPendReg_6 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  excPendReg_7 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  excPendReg_8 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  excPendReg_9 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  excPendReg_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  excPendReg_11 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  excPendReg_12 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  excPendReg_13 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  excPendReg_14 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  excPendReg_15 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  excPendReg_16 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  excPendReg_17 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  excPendReg_18 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  excPendReg_19 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  excPendReg_20 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  excPendReg_21 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  excPendReg_22 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  excPendReg_23 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  excPendReg_24 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  excPendReg_25 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  excPendReg_26 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  excPendReg_27 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  excPendReg_28 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  excPendReg_29 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  excPendReg_30 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  excPendReg_31 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  intrPendReg_16 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  intrPendReg_17 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  intrPendReg_18 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  intrPendReg_19 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  intrPendReg_20 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  intrPendReg_21 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  REG = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  REG_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  REG_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  REG_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  REG_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  REG_5 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  excBaseReg = _RAND_54[29:0];
  _RAND_55 = {1{`RANDOM}};
  excAddrReg = _RAND_55[29:0];
  _RAND_56 = {1{`RANDOM}};
  srcReg = _RAND_56[4:0];
  _RAND_57 = {1{`RANDOM}};
  exc = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  intr = _RAND_58[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemBlock_4(
  input         clock,
  input  [7:0]  io_rdAddr,
  output [19:0] io_rdData,
  input  [7:0]  io_wrAddr,
  input         io_wrEna,
  input  [19:0] io_wrData
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] mem [0:255];
  wire [19:0] mem_MPORT_1_data;
  wire [7:0] mem_MPORT_1_addr;
  wire [19:0] mem_MPORT_data;
  wire [7:0] mem_MPORT_addr;
  wire  mem_MPORT_mask;
  wire  mem_MPORT_en;
  reg [7:0] rdAddrReg; // @[MemBlock.scala 59:22]
  reg  REG; // @[MemBlock.scala 64:14]
  reg [7:0] REG_1; // @[MemBlock.scala 65:14]
  wire  _T_4 = REG_1 == rdAddrReg; // @[MemBlock.scala 65:33]
  wire  _T_5 = REG & _T_4; // @[MemBlock.scala 64:44]
  reg [19:0] REG_2; // @[MemBlock.scala 66:29]
  assign mem_MPORT_1_addr = rdAddrReg;
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr];
  assign mem_MPORT_data = io_wrData;
  assign mem_MPORT_addr = io_wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEna;
  assign io_rdData = _T_5 ? REG_2 : mem_MPORT_1_data; // @[MemBlock.scala 65:48 MemBlock.scala 66:23 MemBlock.scala 60:13]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data;
    end
    rdAddrReg <= io_rdAddr; // @[MemBlock.scala 59:22]
    REG <= io_wrEna; // @[MemBlock.scala 64:14]
    REG_1 <= io_wrAddr; // @[MemBlock.scala 65:14]
    REG_2 <= io_wrData; // @[MemBlock.scala 66:29]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem[initvar] = _RAND_0[19:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rdAddrReg = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_1 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[19:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemBlock_5(
  input        clock,
  input  [9:0] io_rdAddr,
  output [7:0] io_rdData,
  input  [9:0] io_wrAddr,
  input        io_wrEna,
  input  [7:0] io_wrData
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] mem [0:1023];
  wire [7:0] mem_MPORT_1_data;
  wire [9:0] mem_MPORT_1_addr;
  wire [7:0] mem_MPORT_data;
  wire [9:0] mem_MPORT_addr;
  wire  mem_MPORT_mask;
  wire  mem_MPORT_en;
  reg [9:0] rdAddrReg; // @[MemBlock.scala 59:22]
  reg  REG; // @[MemBlock.scala 64:14]
  reg [9:0] REG_1; // @[MemBlock.scala 65:14]
  wire  _T_4 = REG_1 == rdAddrReg; // @[MemBlock.scala 65:33]
  wire  _T_5 = REG & _T_4; // @[MemBlock.scala 64:44]
  reg [7:0] REG_2; // @[MemBlock.scala 66:29]
  assign mem_MPORT_1_addr = rdAddrReg;
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr];
  assign mem_MPORT_data = io_wrData;
  assign mem_MPORT_addr = io_wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEna;
  assign io_rdData = _T_5 ? REG_2 : mem_MPORT_1_data; // @[MemBlock.scala 65:48 MemBlock.scala 66:23 MemBlock.scala 60:13]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data;
    end
    rdAddrReg <= io_rdAddr; // @[MemBlock.scala 59:22]
    REG <= io_wrEna; // @[MemBlock.scala 64:14]
    REG_1 <= io_wrAddr; // @[MemBlock.scala 65:14]
    REG_2 <= io_wrData; // @[MemBlock.scala 66:29]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    mem[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rdAddrReg = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_1 = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DirectMappedCache(
  input         clock,
  input         reset,
  input  [2:0]  io_master_M_Cmd,
  input  [31:0] io_master_M_Addr,
  input  [31:0] io_master_M_Data,
  input  [3:0]  io_master_M_ByteEn,
  output [1:0]  io_master_S_Resp,
  output [31:0] io_master_S_Data,
  output [2:0]  io_slave_M_Cmd,
  output [31:0] io_slave_M_Addr,
  input  [1:0]  io_slave_S_Resp,
  input  [31:0] io_slave_S_Data,
  input         io_slave_S_CmdAccept,
  input         io_invalidate
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
`endif // RANDOMIZE_REG_INIT
  wire  tagMem_clock; // @[MemBlock.scala 15:11]
  wire [7:0] tagMem_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [19:0] tagMem_io_rdData; // @[MemBlock.scala 15:11]
  wire [7:0] tagMem_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  tagMem_io_wrEna; // @[MemBlock.scala 15:11]
  wire [19:0] tagMem_io_wrData; // @[MemBlock.scala 15:11]
  wire  MemBlock_clock; // @[MemBlock.scala 15:11]
  wire [9:0] MemBlock_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_io_rdData; // @[MemBlock.scala 15:11]
  wire [9:0] MemBlock_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_io_wrData; // @[MemBlock.scala 15:11]
  wire  MemBlock_1_clock; // @[MemBlock.scala 15:11]
  wire [9:0] MemBlock_1_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_1_io_rdData; // @[MemBlock.scala 15:11]
  wire [9:0] MemBlock_1_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_1_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_1_io_wrData; // @[MemBlock.scala 15:11]
  wire  MemBlock_2_clock; // @[MemBlock.scala 15:11]
  wire [9:0] MemBlock_2_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_2_io_rdData; // @[MemBlock.scala 15:11]
  wire [9:0] MemBlock_2_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_2_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_2_io_wrData; // @[MemBlock.scala 15:11]
  wire  MemBlock_3_clock; // @[MemBlock.scala 15:11]
  wire [9:0] MemBlock_3_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_3_io_rdData; // @[MemBlock.scala 15:11]
  wire [9:0] MemBlock_3_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_3_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_3_io_wrData; // @[MemBlock.scala 15:11]
  reg [2:0] masterReg_Cmd; // @[DirectMappedCache.scala 37:22]
  reg [31:0] masterReg_Addr; // @[DirectMappedCache.scala 37:22]
  reg [3:0] masterReg_ByteEn; // @[DirectMappedCache.scala 37:22]
  reg  tagVMem_0; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_1; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_2; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_3; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_4; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_5; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_6; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_7; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_8; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_9; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_10; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_11; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_12; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_13; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_14; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_15; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_16; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_17; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_18; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_19; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_20; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_21; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_22; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_23; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_24; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_25; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_26; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_27; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_28; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_29; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_30; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_31; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_32; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_33; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_34; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_35; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_36; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_37; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_38; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_39; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_40; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_41; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_42; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_43; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_44; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_45; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_46; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_47; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_48; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_49; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_50; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_51; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_52; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_53; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_54; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_55; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_56; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_57; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_58; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_59; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_60; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_61; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_62; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_63; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_64; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_65; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_66; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_67; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_68; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_69; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_70; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_71; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_72; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_73; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_74; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_75; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_76; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_77; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_78; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_79; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_80; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_81; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_82; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_83; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_84; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_85; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_86; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_87; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_88; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_89; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_90; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_91; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_92; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_93; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_94; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_95; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_96; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_97; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_98; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_99; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_100; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_101; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_102; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_103; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_104; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_105; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_106; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_107; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_108; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_109; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_110; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_111; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_112; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_113; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_114; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_115; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_116; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_117; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_118; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_119; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_120; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_121; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_122; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_123; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_124; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_125; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_126; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_127; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_128; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_129; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_130; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_131; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_132; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_133; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_134; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_135; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_136; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_137; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_138; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_139; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_140; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_141; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_142; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_143; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_144; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_145; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_146; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_147; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_148; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_149; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_150; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_151; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_152; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_153; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_154; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_155; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_156; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_157; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_158; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_159; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_160; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_161; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_162; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_163; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_164; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_165; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_166; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_167; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_168; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_169; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_170; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_171; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_172; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_173; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_174; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_175; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_176; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_177; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_178; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_179; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_180; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_181; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_182; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_183; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_184; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_185; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_186; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_187; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_188; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_189; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_190; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_191; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_192; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_193; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_194; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_195; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_196; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_197; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_198; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_199; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_200; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_201; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_202; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_203; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_204; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_205; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_206; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_207; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_208; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_209; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_210; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_211; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_212; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_213; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_214; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_215; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_216; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_217; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_218; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_219; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_220; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_221; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_222; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_223; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_224; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_225; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_226; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_227; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_228; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_229; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_230; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_231; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_232; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_233; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_234; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_235; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_236; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_237; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_238; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_239; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_240; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_241; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_242; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_243; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_244; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_245; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_246; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_247; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_248; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_249; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_250; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_251; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_252; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_253; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_254; // @[DirectMappedCache.scala 42:24]
  reg  tagVMem_255; // @[DirectMappedCache.scala 42:24]
  reg  tagV; // @[DirectMappedCache.scala 49:17]
  wire  _GEN_1 = 8'h1 == io_master_M_Addr[11:4] ? tagVMem_1 : tagVMem_0; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_2 = 8'h2 == io_master_M_Addr[11:4] ? tagVMem_2 : _GEN_1; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_3 = 8'h3 == io_master_M_Addr[11:4] ? tagVMem_3 : _GEN_2; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_4 = 8'h4 == io_master_M_Addr[11:4] ? tagVMem_4 : _GEN_3; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_5 = 8'h5 == io_master_M_Addr[11:4] ? tagVMem_5 : _GEN_4; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_6 = 8'h6 == io_master_M_Addr[11:4] ? tagVMem_6 : _GEN_5; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_7 = 8'h7 == io_master_M_Addr[11:4] ? tagVMem_7 : _GEN_6; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_8 = 8'h8 == io_master_M_Addr[11:4] ? tagVMem_8 : _GEN_7; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_9 = 8'h9 == io_master_M_Addr[11:4] ? tagVMem_9 : _GEN_8; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_10 = 8'ha == io_master_M_Addr[11:4] ? tagVMem_10 : _GEN_9; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_11 = 8'hb == io_master_M_Addr[11:4] ? tagVMem_11 : _GEN_10; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_12 = 8'hc == io_master_M_Addr[11:4] ? tagVMem_12 : _GEN_11; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_13 = 8'hd == io_master_M_Addr[11:4] ? tagVMem_13 : _GEN_12; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_14 = 8'he == io_master_M_Addr[11:4] ? tagVMem_14 : _GEN_13; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_15 = 8'hf == io_master_M_Addr[11:4] ? tagVMem_15 : _GEN_14; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_16 = 8'h10 == io_master_M_Addr[11:4] ? tagVMem_16 : _GEN_15; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_17 = 8'h11 == io_master_M_Addr[11:4] ? tagVMem_17 : _GEN_16; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_18 = 8'h12 == io_master_M_Addr[11:4] ? tagVMem_18 : _GEN_17; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_19 = 8'h13 == io_master_M_Addr[11:4] ? tagVMem_19 : _GEN_18; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_20 = 8'h14 == io_master_M_Addr[11:4] ? tagVMem_20 : _GEN_19; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_21 = 8'h15 == io_master_M_Addr[11:4] ? tagVMem_21 : _GEN_20; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_22 = 8'h16 == io_master_M_Addr[11:4] ? tagVMem_22 : _GEN_21; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_23 = 8'h17 == io_master_M_Addr[11:4] ? tagVMem_23 : _GEN_22; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_24 = 8'h18 == io_master_M_Addr[11:4] ? tagVMem_24 : _GEN_23; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_25 = 8'h19 == io_master_M_Addr[11:4] ? tagVMem_25 : _GEN_24; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_26 = 8'h1a == io_master_M_Addr[11:4] ? tagVMem_26 : _GEN_25; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_27 = 8'h1b == io_master_M_Addr[11:4] ? tagVMem_27 : _GEN_26; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_28 = 8'h1c == io_master_M_Addr[11:4] ? tagVMem_28 : _GEN_27; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_29 = 8'h1d == io_master_M_Addr[11:4] ? tagVMem_29 : _GEN_28; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_30 = 8'h1e == io_master_M_Addr[11:4] ? tagVMem_30 : _GEN_29; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_31 = 8'h1f == io_master_M_Addr[11:4] ? tagVMem_31 : _GEN_30; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_32 = 8'h20 == io_master_M_Addr[11:4] ? tagVMem_32 : _GEN_31; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_33 = 8'h21 == io_master_M_Addr[11:4] ? tagVMem_33 : _GEN_32; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_34 = 8'h22 == io_master_M_Addr[11:4] ? tagVMem_34 : _GEN_33; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_35 = 8'h23 == io_master_M_Addr[11:4] ? tagVMem_35 : _GEN_34; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_36 = 8'h24 == io_master_M_Addr[11:4] ? tagVMem_36 : _GEN_35; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_37 = 8'h25 == io_master_M_Addr[11:4] ? tagVMem_37 : _GEN_36; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_38 = 8'h26 == io_master_M_Addr[11:4] ? tagVMem_38 : _GEN_37; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_39 = 8'h27 == io_master_M_Addr[11:4] ? tagVMem_39 : _GEN_38; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_40 = 8'h28 == io_master_M_Addr[11:4] ? tagVMem_40 : _GEN_39; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_41 = 8'h29 == io_master_M_Addr[11:4] ? tagVMem_41 : _GEN_40; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_42 = 8'h2a == io_master_M_Addr[11:4] ? tagVMem_42 : _GEN_41; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_43 = 8'h2b == io_master_M_Addr[11:4] ? tagVMem_43 : _GEN_42; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_44 = 8'h2c == io_master_M_Addr[11:4] ? tagVMem_44 : _GEN_43; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_45 = 8'h2d == io_master_M_Addr[11:4] ? tagVMem_45 : _GEN_44; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_46 = 8'h2e == io_master_M_Addr[11:4] ? tagVMem_46 : _GEN_45; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_47 = 8'h2f == io_master_M_Addr[11:4] ? tagVMem_47 : _GEN_46; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_48 = 8'h30 == io_master_M_Addr[11:4] ? tagVMem_48 : _GEN_47; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_49 = 8'h31 == io_master_M_Addr[11:4] ? tagVMem_49 : _GEN_48; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_50 = 8'h32 == io_master_M_Addr[11:4] ? tagVMem_50 : _GEN_49; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_51 = 8'h33 == io_master_M_Addr[11:4] ? tagVMem_51 : _GEN_50; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_52 = 8'h34 == io_master_M_Addr[11:4] ? tagVMem_52 : _GEN_51; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_53 = 8'h35 == io_master_M_Addr[11:4] ? tagVMem_53 : _GEN_52; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_54 = 8'h36 == io_master_M_Addr[11:4] ? tagVMem_54 : _GEN_53; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_55 = 8'h37 == io_master_M_Addr[11:4] ? tagVMem_55 : _GEN_54; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_56 = 8'h38 == io_master_M_Addr[11:4] ? tagVMem_56 : _GEN_55; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_57 = 8'h39 == io_master_M_Addr[11:4] ? tagVMem_57 : _GEN_56; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_58 = 8'h3a == io_master_M_Addr[11:4] ? tagVMem_58 : _GEN_57; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_59 = 8'h3b == io_master_M_Addr[11:4] ? tagVMem_59 : _GEN_58; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_60 = 8'h3c == io_master_M_Addr[11:4] ? tagVMem_60 : _GEN_59; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_61 = 8'h3d == io_master_M_Addr[11:4] ? tagVMem_61 : _GEN_60; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_62 = 8'h3e == io_master_M_Addr[11:4] ? tagVMem_62 : _GEN_61; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_63 = 8'h3f == io_master_M_Addr[11:4] ? tagVMem_63 : _GEN_62; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_64 = 8'h40 == io_master_M_Addr[11:4] ? tagVMem_64 : _GEN_63; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_65 = 8'h41 == io_master_M_Addr[11:4] ? tagVMem_65 : _GEN_64; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_66 = 8'h42 == io_master_M_Addr[11:4] ? tagVMem_66 : _GEN_65; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_67 = 8'h43 == io_master_M_Addr[11:4] ? tagVMem_67 : _GEN_66; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_68 = 8'h44 == io_master_M_Addr[11:4] ? tagVMem_68 : _GEN_67; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_69 = 8'h45 == io_master_M_Addr[11:4] ? tagVMem_69 : _GEN_68; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_70 = 8'h46 == io_master_M_Addr[11:4] ? tagVMem_70 : _GEN_69; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_71 = 8'h47 == io_master_M_Addr[11:4] ? tagVMem_71 : _GEN_70; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_72 = 8'h48 == io_master_M_Addr[11:4] ? tagVMem_72 : _GEN_71; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_73 = 8'h49 == io_master_M_Addr[11:4] ? tagVMem_73 : _GEN_72; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_74 = 8'h4a == io_master_M_Addr[11:4] ? tagVMem_74 : _GEN_73; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_75 = 8'h4b == io_master_M_Addr[11:4] ? tagVMem_75 : _GEN_74; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_76 = 8'h4c == io_master_M_Addr[11:4] ? tagVMem_76 : _GEN_75; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_77 = 8'h4d == io_master_M_Addr[11:4] ? tagVMem_77 : _GEN_76; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_78 = 8'h4e == io_master_M_Addr[11:4] ? tagVMem_78 : _GEN_77; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_79 = 8'h4f == io_master_M_Addr[11:4] ? tagVMem_79 : _GEN_78; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_80 = 8'h50 == io_master_M_Addr[11:4] ? tagVMem_80 : _GEN_79; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_81 = 8'h51 == io_master_M_Addr[11:4] ? tagVMem_81 : _GEN_80; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_82 = 8'h52 == io_master_M_Addr[11:4] ? tagVMem_82 : _GEN_81; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_83 = 8'h53 == io_master_M_Addr[11:4] ? tagVMem_83 : _GEN_82; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_84 = 8'h54 == io_master_M_Addr[11:4] ? tagVMem_84 : _GEN_83; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_85 = 8'h55 == io_master_M_Addr[11:4] ? tagVMem_85 : _GEN_84; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_86 = 8'h56 == io_master_M_Addr[11:4] ? tagVMem_86 : _GEN_85; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_87 = 8'h57 == io_master_M_Addr[11:4] ? tagVMem_87 : _GEN_86; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_88 = 8'h58 == io_master_M_Addr[11:4] ? tagVMem_88 : _GEN_87; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_89 = 8'h59 == io_master_M_Addr[11:4] ? tagVMem_89 : _GEN_88; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_90 = 8'h5a == io_master_M_Addr[11:4] ? tagVMem_90 : _GEN_89; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_91 = 8'h5b == io_master_M_Addr[11:4] ? tagVMem_91 : _GEN_90; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_92 = 8'h5c == io_master_M_Addr[11:4] ? tagVMem_92 : _GEN_91; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_93 = 8'h5d == io_master_M_Addr[11:4] ? tagVMem_93 : _GEN_92; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_94 = 8'h5e == io_master_M_Addr[11:4] ? tagVMem_94 : _GEN_93; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_95 = 8'h5f == io_master_M_Addr[11:4] ? tagVMem_95 : _GEN_94; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_96 = 8'h60 == io_master_M_Addr[11:4] ? tagVMem_96 : _GEN_95; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_97 = 8'h61 == io_master_M_Addr[11:4] ? tagVMem_97 : _GEN_96; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_98 = 8'h62 == io_master_M_Addr[11:4] ? tagVMem_98 : _GEN_97; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_99 = 8'h63 == io_master_M_Addr[11:4] ? tagVMem_99 : _GEN_98; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_100 = 8'h64 == io_master_M_Addr[11:4] ? tagVMem_100 : _GEN_99; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_101 = 8'h65 == io_master_M_Addr[11:4] ? tagVMem_101 : _GEN_100; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_102 = 8'h66 == io_master_M_Addr[11:4] ? tagVMem_102 : _GEN_101; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_103 = 8'h67 == io_master_M_Addr[11:4] ? tagVMem_103 : _GEN_102; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_104 = 8'h68 == io_master_M_Addr[11:4] ? tagVMem_104 : _GEN_103; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_105 = 8'h69 == io_master_M_Addr[11:4] ? tagVMem_105 : _GEN_104; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_106 = 8'h6a == io_master_M_Addr[11:4] ? tagVMem_106 : _GEN_105; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_107 = 8'h6b == io_master_M_Addr[11:4] ? tagVMem_107 : _GEN_106; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_108 = 8'h6c == io_master_M_Addr[11:4] ? tagVMem_108 : _GEN_107; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_109 = 8'h6d == io_master_M_Addr[11:4] ? tagVMem_109 : _GEN_108; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_110 = 8'h6e == io_master_M_Addr[11:4] ? tagVMem_110 : _GEN_109; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_111 = 8'h6f == io_master_M_Addr[11:4] ? tagVMem_111 : _GEN_110; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_112 = 8'h70 == io_master_M_Addr[11:4] ? tagVMem_112 : _GEN_111; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_113 = 8'h71 == io_master_M_Addr[11:4] ? tagVMem_113 : _GEN_112; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_114 = 8'h72 == io_master_M_Addr[11:4] ? tagVMem_114 : _GEN_113; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_115 = 8'h73 == io_master_M_Addr[11:4] ? tagVMem_115 : _GEN_114; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_116 = 8'h74 == io_master_M_Addr[11:4] ? tagVMem_116 : _GEN_115; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_117 = 8'h75 == io_master_M_Addr[11:4] ? tagVMem_117 : _GEN_116; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_118 = 8'h76 == io_master_M_Addr[11:4] ? tagVMem_118 : _GEN_117; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_119 = 8'h77 == io_master_M_Addr[11:4] ? tagVMem_119 : _GEN_118; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_120 = 8'h78 == io_master_M_Addr[11:4] ? tagVMem_120 : _GEN_119; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_121 = 8'h79 == io_master_M_Addr[11:4] ? tagVMem_121 : _GEN_120; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_122 = 8'h7a == io_master_M_Addr[11:4] ? tagVMem_122 : _GEN_121; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_123 = 8'h7b == io_master_M_Addr[11:4] ? tagVMem_123 : _GEN_122; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_124 = 8'h7c == io_master_M_Addr[11:4] ? tagVMem_124 : _GEN_123; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_125 = 8'h7d == io_master_M_Addr[11:4] ? tagVMem_125 : _GEN_124; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_126 = 8'h7e == io_master_M_Addr[11:4] ? tagVMem_126 : _GEN_125; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_127 = 8'h7f == io_master_M_Addr[11:4] ? tagVMem_127 : _GEN_126; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_128 = 8'h80 == io_master_M_Addr[11:4] ? tagVMem_128 : _GEN_127; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_129 = 8'h81 == io_master_M_Addr[11:4] ? tagVMem_129 : _GEN_128; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_130 = 8'h82 == io_master_M_Addr[11:4] ? tagVMem_130 : _GEN_129; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_131 = 8'h83 == io_master_M_Addr[11:4] ? tagVMem_131 : _GEN_130; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_132 = 8'h84 == io_master_M_Addr[11:4] ? tagVMem_132 : _GEN_131; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_133 = 8'h85 == io_master_M_Addr[11:4] ? tagVMem_133 : _GEN_132; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_134 = 8'h86 == io_master_M_Addr[11:4] ? tagVMem_134 : _GEN_133; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_135 = 8'h87 == io_master_M_Addr[11:4] ? tagVMem_135 : _GEN_134; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_136 = 8'h88 == io_master_M_Addr[11:4] ? tagVMem_136 : _GEN_135; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_137 = 8'h89 == io_master_M_Addr[11:4] ? tagVMem_137 : _GEN_136; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_138 = 8'h8a == io_master_M_Addr[11:4] ? tagVMem_138 : _GEN_137; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_139 = 8'h8b == io_master_M_Addr[11:4] ? tagVMem_139 : _GEN_138; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_140 = 8'h8c == io_master_M_Addr[11:4] ? tagVMem_140 : _GEN_139; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_141 = 8'h8d == io_master_M_Addr[11:4] ? tagVMem_141 : _GEN_140; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_142 = 8'h8e == io_master_M_Addr[11:4] ? tagVMem_142 : _GEN_141; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_143 = 8'h8f == io_master_M_Addr[11:4] ? tagVMem_143 : _GEN_142; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_144 = 8'h90 == io_master_M_Addr[11:4] ? tagVMem_144 : _GEN_143; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_145 = 8'h91 == io_master_M_Addr[11:4] ? tagVMem_145 : _GEN_144; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_146 = 8'h92 == io_master_M_Addr[11:4] ? tagVMem_146 : _GEN_145; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_147 = 8'h93 == io_master_M_Addr[11:4] ? tagVMem_147 : _GEN_146; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_148 = 8'h94 == io_master_M_Addr[11:4] ? tagVMem_148 : _GEN_147; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_149 = 8'h95 == io_master_M_Addr[11:4] ? tagVMem_149 : _GEN_148; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_150 = 8'h96 == io_master_M_Addr[11:4] ? tagVMem_150 : _GEN_149; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_151 = 8'h97 == io_master_M_Addr[11:4] ? tagVMem_151 : _GEN_150; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_152 = 8'h98 == io_master_M_Addr[11:4] ? tagVMem_152 : _GEN_151; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_153 = 8'h99 == io_master_M_Addr[11:4] ? tagVMem_153 : _GEN_152; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_154 = 8'h9a == io_master_M_Addr[11:4] ? tagVMem_154 : _GEN_153; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_155 = 8'h9b == io_master_M_Addr[11:4] ? tagVMem_155 : _GEN_154; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_156 = 8'h9c == io_master_M_Addr[11:4] ? tagVMem_156 : _GEN_155; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_157 = 8'h9d == io_master_M_Addr[11:4] ? tagVMem_157 : _GEN_156; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_158 = 8'h9e == io_master_M_Addr[11:4] ? tagVMem_158 : _GEN_157; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_159 = 8'h9f == io_master_M_Addr[11:4] ? tagVMem_159 : _GEN_158; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_160 = 8'ha0 == io_master_M_Addr[11:4] ? tagVMem_160 : _GEN_159; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_161 = 8'ha1 == io_master_M_Addr[11:4] ? tagVMem_161 : _GEN_160; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_162 = 8'ha2 == io_master_M_Addr[11:4] ? tagVMem_162 : _GEN_161; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_163 = 8'ha3 == io_master_M_Addr[11:4] ? tagVMem_163 : _GEN_162; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_164 = 8'ha4 == io_master_M_Addr[11:4] ? tagVMem_164 : _GEN_163; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_165 = 8'ha5 == io_master_M_Addr[11:4] ? tagVMem_165 : _GEN_164; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_166 = 8'ha6 == io_master_M_Addr[11:4] ? tagVMem_166 : _GEN_165; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_167 = 8'ha7 == io_master_M_Addr[11:4] ? tagVMem_167 : _GEN_166; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_168 = 8'ha8 == io_master_M_Addr[11:4] ? tagVMem_168 : _GEN_167; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_169 = 8'ha9 == io_master_M_Addr[11:4] ? tagVMem_169 : _GEN_168; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_170 = 8'haa == io_master_M_Addr[11:4] ? tagVMem_170 : _GEN_169; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_171 = 8'hab == io_master_M_Addr[11:4] ? tagVMem_171 : _GEN_170; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_172 = 8'hac == io_master_M_Addr[11:4] ? tagVMem_172 : _GEN_171; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_173 = 8'had == io_master_M_Addr[11:4] ? tagVMem_173 : _GEN_172; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_174 = 8'hae == io_master_M_Addr[11:4] ? tagVMem_174 : _GEN_173; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_175 = 8'haf == io_master_M_Addr[11:4] ? tagVMem_175 : _GEN_174; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_176 = 8'hb0 == io_master_M_Addr[11:4] ? tagVMem_176 : _GEN_175; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_177 = 8'hb1 == io_master_M_Addr[11:4] ? tagVMem_177 : _GEN_176; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_178 = 8'hb2 == io_master_M_Addr[11:4] ? tagVMem_178 : _GEN_177; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_179 = 8'hb3 == io_master_M_Addr[11:4] ? tagVMem_179 : _GEN_178; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_180 = 8'hb4 == io_master_M_Addr[11:4] ? tagVMem_180 : _GEN_179; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_181 = 8'hb5 == io_master_M_Addr[11:4] ? tagVMem_181 : _GEN_180; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_182 = 8'hb6 == io_master_M_Addr[11:4] ? tagVMem_182 : _GEN_181; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_183 = 8'hb7 == io_master_M_Addr[11:4] ? tagVMem_183 : _GEN_182; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_184 = 8'hb8 == io_master_M_Addr[11:4] ? tagVMem_184 : _GEN_183; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_185 = 8'hb9 == io_master_M_Addr[11:4] ? tagVMem_185 : _GEN_184; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_186 = 8'hba == io_master_M_Addr[11:4] ? tagVMem_186 : _GEN_185; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_187 = 8'hbb == io_master_M_Addr[11:4] ? tagVMem_187 : _GEN_186; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_188 = 8'hbc == io_master_M_Addr[11:4] ? tagVMem_188 : _GEN_187; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_189 = 8'hbd == io_master_M_Addr[11:4] ? tagVMem_189 : _GEN_188; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_190 = 8'hbe == io_master_M_Addr[11:4] ? tagVMem_190 : _GEN_189; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_191 = 8'hbf == io_master_M_Addr[11:4] ? tagVMem_191 : _GEN_190; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_192 = 8'hc0 == io_master_M_Addr[11:4] ? tagVMem_192 : _GEN_191; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_193 = 8'hc1 == io_master_M_Addr[11:4] ? tagVMem_193 : _GEN_192; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_194 = 8'hc2 == io_master_M_Addr[11:4] ? tagVMem_194 : _GEN_193; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_195 = 8'hc3 == io_master_M_Addr[11:4] ? tagVMem_195 : _GEN_194; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_196 = 8'hc4 == io_master_M_Addr[11:4] ? tagVMem_196 : _GEN_195; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_197 = 8'hc5 == io_master_M_Addr[11:4] ? tagVMem_197 : _GEN_196; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_198 = 8'hc6 == io_master_M_Addr[11:4] ? tagVMem_198 : _GEN_197; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_199 = 8'hc7 == io_master_M_Addr[11:4] ? tagVMem_199 : _GEN_198; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_200 = 8'hc8 == io_master_M_Addr[11:4] ? tagVMem_200 : _GEN_199; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_201 = 8'hc9 == io_master_M_Addr[11:4] ? tagVMem_201 : _GEN_200; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_202 = 8'hca == io_master_M_Addr[11:4] ? tagVMem_202 : _GEN_201; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_203 = 8'hcb == io_master_M_Addr[11:4] ? tagVMem_203 : _GEN_202; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_204 = 8'hcc == io_master_M_Addr[11:4] ? tagVMem_204 : _GEN_203; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_205 = 8'hcd == io_master_M_Addr[11:4] ? tagVMem_205 : _GEN_204; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_206 = 8'hce == io_master_M_Addr[11:4] ? tagVMem_206 : _GEN_205; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_207 = 8'hcf == io_master_M_Addr[11:4] ? tagVMem_207 : _GEN_206; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_208 = 8'hd0 == io_master_M_Addr[11:4] ? tagVMem_208 : _GEN_207; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_209 = 8'hd1 == io_master_M_Addr[11:4] ? tagVMem_209 : _GEN_208; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_210 = 8'hd2 == io_master_M_Addr[11:4] ? tagVMem_210 : _GEN_209; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_211 = 8'hd3 == io_master_M_Addr[11:4] ? tagVMem_211 : _GEN_210; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_212 = 8'hd4 == io_master_M_Addr[11:4] ? tagVMem_212 : _GEN_211; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_213 = 8'hd5 == io_master_M_Addr[11:4] ? tagVMem_213 : _GEN_212; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_214 = 8'hd6 == io_master_M_Addr[11:4] ? tagVMem_214 : _GEN_213; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_215 = 8'hd7 == io_master_M_Addr[11:4] ? tagVMem_215 : _GEN_214; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_216 = 8'hd8 == io_master_M_Addr[11:4] ? tagVMem_216 : _GEN_215; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_217 = 8'hd9 == io_master_M_Addr[11:4] ? tagVMem_217 : _GEN_216; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_218 = 8'hda == io_master_M_Addr[11:4] ? tagVMem_218 : _GEN_217; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_219 = 8'hdb == io_master_M_Addr[11:4] ? tagVMem_219 : _GEN_218; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_220 = 8'hdc == io_master_M_Addr[11:4] ? tagVMem_220 : _GEN_219; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_221 = 8'hdd == io_master_M_Addr[11:4] ? tagVMem_221 : _GEN_220; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_222 = 8'hde == io_master_M_Addr[11:4] ? tagVMem_222 : _GEN_221; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_223 = 8'hdf == io_master_M_Addr[11:4] ? tagVMem_223 : _GEN_222; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_224 = 8'he0 == io_master_M_Addr[11:4] ? tagVMem_224 : _GEN_223; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_225 = 8'he1 == io_master_M_Addr[11:4] ? tagVMem_225 : _GEN_224; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_226 = 8'he2 == io_master_M_Addr[11:4] ? tagVMem_226 : _GEN_225; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_227 = 8'he3 == io_master_M_Addr[11:4] ? tagVMem_227 : _GEN_226; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_228 = 8'he4 == io_master_M_Addr[11:4] ? tagVMem_228 : _GEN_227; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_229 = 8'he5 == io_master_M_Addr[11:4] ? tagVMem_229 : _GEN_228; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_230 = 8'he6 == io_master_M_Addr[11:4] ? tagVMem_230 : _GEN_229; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_231 = 8'he7 == io_master_M_Addr[11:4] ? tagVMem_231 : _GEN_230; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_232 = 8'he8 == io_master_M_Addr[11:4] ? tagVMem_232 : _GEN_231; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_233 = 8'he9 == io_master_M_Addr[11:4] ? tagVMem_233 : _GEN_232; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_234 = 8'hea == io_master_M_Addr[11:4] ? tagVMem_234 : _GEN_233; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_235 = 8'heb == io_master_M_Addr[11:4] ? tagVMem_235 : _GEN_234; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_236 = 8'hec == io_master_M_Addr[11:4] ? tagVMem_236 : _GEN_235; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_237 = 8'hed == io_master_M_Addr[11:4] ? tagVMem_237 : _GEN_236; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_238 = 8'hee == io_master_M_Addr[11:4] ? tagVMem_238 : _GEN_237; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_239 = 8'hef == io_master_M_Addr[11:4] ? tagVMem_239 : _GEN_238; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_240 = 8'hf0 == io_master_M_Addr[11:4] ? tagVMem_240 : _GEN_239; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_241 = 8'hf1 == io_master_M_Addr[11:4] ? tagVMem_241 : _GEN_240; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_242 = 8'hf2 == io_master_M_Addr[11:4] ? tagVMem_242 : _GEN_241; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_243 = 8'hf3 == io_master_M_Addr[11:4] ? tagVMem_243 : _GEN_242; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_244 = 8'hf4 == io_master_M_Addr[11:4] ? tagVMem_244 : _GEN_243; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_245 = 8'hf5 == io_master_M_Addr[11:4] ? tagVMem_245 : _GEN_244; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_246 = 8'hf6 == io_master_M_Addr[11:4] ? tagVMem_246 : _GEN_245; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_247 = 8'hf7 == io_master_M_Addr[11:4] ? tagVMem_247 : _GEN_246; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_248 = 8'hf8 == io_master_M_Addr[11:4] ? tagVMem_248 : _GEN_247; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_249 = 8'hf9 == io_master_M_Addr[11:4] ? tagVMem_249 : _GEN_248; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_250 = 8'hfa == io_master_M_Addr[11:4] ? tagVMem_250 : _GEN_249; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  _GEN_251 = 8'hfb == io_master_M_Addr[11:4] ? tagVMem_251 : _GEN_250; // @[DirectMappedCache.scala 49:17 DirectMappedCache.scala 49:17]
  wire  tagValid = tagV & tagMem_io_rdData == masterReg_Addr[31:12]; // @[DirectMappedCache.scala 50:23]
  reg  fillReg; // @[DirectMappedCache.scala 52:20]
  reg [9:0] wrAddrReg; // @[DirectMappedCache.scala 54:22]
  reg [31:0] wrDataReg; // @[DirectMappedCache.scala 55:22]
  wire [3:0] stmsk = masterReg_Cmd == 3'h1 ? masterReg_ByteEn : 4'h0; // @[DirectMappedCache.scala 61:18]
  wire [31:0] rdData = {MemBlock_3_io_rdData,MemBlock_2_io_rdData,MemBlock_1_io_rdData,MemBlock_io_rdData}; // @[DirectMappedCache.scala 68:84]
  wire  _T_28 = masterReg_Cmd == 3'h2; // @[DirectMappedCache.scala 72:53]
  wire [1:0] _T_30 = tagValid & masterReg_Cmd == 3'h2 ? 2'h1 : 2'h0; // @[DirectMappedCache.scala 72:26]
  reg [1:0] stateReg; // @[DirectMappedCache.scala 77:21]
  reg [1:0] burstCntReg; // @[DirectMappedCache.scala 79:24]
  reg [1:0] missIndexReg; // @[DirectMappedCache.scala 80:25]
  reg [1:0] slaveReg_Resp; // @[DirectMappedCache.scala 83:21]
  reg [31:0] slaveReg_Data; // @[DirectMappedCache.scala 83:21]
  wire [27:0] hi = masterReg_Addr[31:4]; // @[DirectMappedCache.scala 87:40]
  wire  _T_34 = ~tagValid; // @[DirectMappedCache.scala 101:8]
  wire  _GEN_257 = 8'h0 == masterReg_Addr[11:4] | tagVMem_0; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_258 = 8'h1 == masterReg_Addr[11:4] | tagVMem_1; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_259 = 8'h2 == masterReg_Addr[11:4] | tagVMem_2; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_260 = 8'h3 == masterReg_Addr[11:4] | tagVMem_3; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_261 = 8'h4 == masterReg_Addr[11:4] | tagVMem_4; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_262 = 8'h5 == masterReg_Addr[11:4] | tagVMem_5; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_263 = 8'h6 == masterReg_Addr[11:4] | tagVMem_6; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_264 = 8'h7 == masterReg_Addr[11:4] | tagVMem_7; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_265 = 8'h8 == masterReg_Addr[11:4] | tagVMem_8; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_266 = 8'h9 == masterReg_Addr[11:4] | tagVMem_9; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_267 = 8'ha == masterReg_Addr[11:4] | tagVMem_10; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_268 = 8'hb == masterReg_Addr[11:4] | tagVMem_11; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_269 = 8'hc == masterReg_Addr[11:4] | tagVMem_12; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_270 = 8'hd == masterReg_Addr[11:4] | tagVMem_13; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_271 = 8'he == masterReg_Addr[11:4] | tagVMem_14; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_272 = 8'hf == masterReg_Addr[11:4] | tagVMem_15; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_273 = 8'h10 == masterReg_Addr[11:4] | tagVMem_16; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_274 = 8'h11 == masterReg_Addr[11:4] | tagVMem_17; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_275 = 8'h12 == masterReg_Addr[11:4] | tagVMem_18; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_276 = 8'h13 == masterReg_Addr[11:4] | tagVMem_19; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_277 = 8'h14 == masterReg_Addr[11:4] | tagVMem_20; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_278 = 8'h15 == masterReg_Addr[11:4] | tagVMem_21; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_279 = 8'h16 == masterReg_Addr[11:4] | tagVMem_22; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_280 = 8'h17 == masterReg_Addr[11:4] | tagVMem_23; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_281 = 8'h18 == masterReg_Addr[11:4] | tagVMem_24; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_282 = 8'h19 == masterReg_Addr[11:4] | tagVMem_25; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_283 = 8'h1a == masterReg_Addr[11:4] | tagVMem_26; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_284 = 8'h1b == masterReg_Addr[11:4] | tagVMem_27; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_285 = 8'h1c == masterReg_Addr[11:4] | tagVMem_28; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_286 = 8'h1d == masterReg_Addr[11:4] | tagVMem_29; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_287 = 8'h1e == masterReg_Addr[11:4] | tagVMem_30; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_288 = 8'h1f == masterReg_Addr[11:4] | tagVMem_31; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_289 = 8'h20 == masterReg_Addr[11:4] | tagVMem_32; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_290 = 8'h21 == masterReg_Addr[11:4] | tagVMem_33; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_291 = 8'h22 == masterReg_Addr[11:4] | tagVMem_34; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_292 = 8'h23 == masterReg_Addr[11:4] | tagVMem_35; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_293 = 8'h24 == masterReg_Addr[11:4] | tagVMem_36; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_294 = 8'h25 == masterReg_Addr[11:4] | tagVMem_37; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_295 = 8'h26 == masterReg_Addr[11:4] | tagVMem_38; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_296 = 8'h27 == masterReg_Addr[11:4] | tagVMem_39; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_297 = 8'h28 == masterReg_Addr[11:4] | tagVMem_40; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_298 = 8'h29 == masterReg_Addr[11:4] | tagVMem_41; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_299 = 8'h2a == masterReg_Addr[11:4] | tagVMem_42; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_300 = 8'h2b == masterReg_Addr[11:4] | tagVMem_43; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_301 = 8'h2c == masterReg_Addr[11:4] | tagVMem_44; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_302 = 8'h2d == masterReg_Addr[11:4] | tagVMem_45; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_303 = 8'h2e == masterReg_Addr[11:4] | tagVMem_46; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_304 = 8'h2f == masterReg_Addr[11:4] | tagVMem_47; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_305 = 8'h30 == masterReg_Addr[11:4] | tagVMem_48; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_306 = 8'h31 == masterReg_Addr[11:4] | tagVMem_49; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_307 = 8'h32 == masterReg_Addr[11:4] | tagVMem_50; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_308 = 8'h33 == masterReg_Addr[11:4] | tagVMem_51; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_309 = 8'h34 == masterReg_Addr[11:4] | tagVMem_52; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_310 = 8'h35 == masterReg_Addr[11:4] | tagVMem_53; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_311 = 8'h36 == masterReg_Addr[11:4] | tagVMem_54; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_312 = 8'h37 == masterReg_Addr[11:4] | tagVMem_55; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_313 = 8'h38 == masterReg_Addr[11:4] | tagVMem_56; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_314 = 8'h39 == masterReg_Addr[11:4] | tagVMem_57; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_315 = 8'h3a == masterReg_Addr[11:4] | tagVMem_58; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_316 = 8'h3b == masterReg_Addr[11:4] | tagVMem_59; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_317 = 8'h3c == masterReg_Addr[11:4] | tagVMem_60; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_318 = 8'h3d == masterReg_Addr[11:4] | tagVMem_61; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_319 = 8'h3e == masterReg_Addr[11:4] | tagVMem_62; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_320 = 8'h3f == masterReg_Addr[11:4] | tagVMem_63; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_321 = 8'h40 == masterReg_Addr[11:4] | tagVMem_64; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_322 = 8'h41 == masterReg_Addr[11:4] | tagVMem_65; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_323 = 8'h42 == masterReg_Addr[11:4] | tagVMem_66; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_324 = 8'h43 == masterReg_Addr[11:4] | tagVMem_67; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_325 = 8'h44 == masterReg_Addr[11:4] | tagVMem_68; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_326 = 8'h45 == masterReg_Addr[11:4] | tagVMem_69; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_327 = 8'h46 == masterReg_Addr[11:4] | tagVMem_70; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_328 = 8'h47 == masterReg_Addr[11:4] | tagVMem_71; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_329 = 8'h48 == masterReg_Addr[11:4] | tagVMem_72; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_330 = 8'h49 == masterReg_Addr[11:4] | tagVMem_73; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_331 = 8'h4a == masterReg_Addr[11:4] | tagVMem_74; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_332 = 8'h4b == masterReg_Addr[11:4] | tagVMem_75; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_333 = 8'h4c == masterReg_Addr[11:4] | tagVMem_76; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_334 = 8'h4d == masterReg_Addr[11:4] | tagVMem_77; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_335 = 8'h4e == masterReg_Addr[11:4] | tagVMem_78; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_336 = 8'h4f == masterReg_Addr[11:4] | tagVMem_79; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_337 = 8'h50 == masterReg_Addr[11:4] | tagVMem_80; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_338 = 8'h51 == masterReg_Addr[11:4] | tagVMem_81; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_339 = 8'h52 == masterReg_Addr[11:4] | tagVMem_82; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_340 = 8'h53 == masterReg_Addr[11:4] | tagVMem_83; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_341 = 8'h54 == masterReg_Addr[11:4] | tagVMem_84; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_342 = 8'h55 == masterReg_Addr[11:4] | tagVMem_85; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_343 = 8'h56 == masterReg_Addr[11:4] | tagVMem_86; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_344 = 8'h57 == masterReg_Addr[11:4] | tagVMem_87; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_345 = 8'h58 == masterReg_Addr[11:4] | tagVMem_88; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_346 = 8'h59 == masterReg_Addr[11:4] | tagVMem_89; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_347 = 8'h5a == masterReg_Addr[11:4] | tagVMem_90; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_348 = 8'h5b == masterReg_Addr[11:4] | tagVMem_91; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_349 = 8'h5c == masterReg_Addr[11:4] | tagVMem_92; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_350 = 8'h5d == masterReg_Addr[11:4] | tagVMem_93; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_351 = 8'h5e == masterReg_Addr[11:4] | tagVMem_94; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_352 = 8'h5f == masterReg_Addr[11:4] | tagVMem_95; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_353 = 8'h60 == masterReg_Addr[11:4] | tagVMem_96; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_354 = 8'h61 == masterReg_Addr[11:4] | tagVMem_97; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_355 = 8'h62 == masterReg_Addr[11:4] | tagVMem_98; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_356 = 8'h63 == masterReg_Addr[11:4] | tagVMem_99; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_357 = 8'h64 == masterReg_Addr[11:4] | tagVMem_100; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_358 = 8'h65 == masterReg_Addr[11:4] | tagVMem_101; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_359 = 8'h66 == masterReg_Addr[11:4] | tagVMem_102; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_360 = 8'h67 == masterReg_Addr[11:4] | tagVMem_103; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_361 = 8'h68 == masterReg_Addr[11:4] | tagVMem_104; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_362 = 8'h69 == masterReg_Addr[11:4] | tagVMem_105; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_363 = 8'h6a == masterReg_Addr[11:4] | tagVMem_106; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_364 = 8'h6b == masterReg_Addr[11:4] | tagVMem_107; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_365 = 8'h6c == masterReg_Addr[11:4] | tagVMem_108; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_366 = 8'h6d == masterReg_Addr[11:4] | tagVMem_109; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_367 = 8'h6e == masterReg_Addr[11:4] | tagVMem_110; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_368 = 8'h6f == masterReg_Addr[11:4] | tagVMem_111; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_369 = 8'h70 == masterReg_Addr[11:4] | tagVMem_112; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_370 = 8'h71 == masterReg_Addr[11:4] | tagVMem_113; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_371 = 8'h72 == masterReg_Addr[11:4] | tagVMem_114; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_372 = 8'h73 == masterReg_Addr[11:4] | tagVMem_115; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_373 = 8'h74 == masterReg_Addr[11:4] | tagVMem_116; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_374 = 8'h75 == masterReg_Addr[11:4] | tagVMem_117; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_375 = 8'h76 == masterReg_Addr[11:4] | tagVMem_118; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_376 = 8'h77 == masterReg_Addr[11:4] | tagVMem_119; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_377 = 8'h78 == masterReg_Addr[11:4] | tagVMem_120; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_378 = 8'h79 == masterReg_Addr[11:4] | tagVMem_121; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_379 = 8'h7a == masterReg_Addr[11:4] | tagVMem_122; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_380 = 8'h7b == masterReg_Addr[11:4] | tagVMem_123; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_381 = 8'h7c == masterReg_Addr[11:4] | tagVMem_124; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_382 = 8'h7d == masterReg_Addr[11:4] | tagVMem_125; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_383 = 8'h7e == masterReg_Addr[11:4] | tagVMem_126; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_384 = 8'h7f == masterReg_Addr[11:4] | tagVMem_127; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_385 = 8'h80 == masterReg_Addr[11:4] | tagVMem_128; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_386 = 8'h81 == masterReg_Addr[11:4] | tagVMem_129; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_387 = 8'h82 == masterReg_Addr[11:4] | tagVMem_130; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_388 = 8'h83 == masterReg_Addr[11:4] | tagVMem_131; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_389 = 8'h84 == masterReg_Addr[11:4] | tagVMem_132; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_390 = 8'h85 == masterReg_Addr[11:4] | tagVMem_133; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_391 = 8'h86 == masterReg_Addr[11:4] | tagVMem_134; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_392 = 8'h87 == masterReg_Addr[11:4] | tagVMem_135; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_393 = 8'h88 == masterReg_Addr[11:4] | tagVMem_136; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_394 = 8'h89 == masterReg_Addr[11:4] | tagVMem_137; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_395 = 8'h8a == masterReg_Addr[11:4] | tagVMem_138; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_396 = 8'h8b == masterReg_Addr[11:4] | tagVMem_139; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_397 = 8'h8c == masterReg_Addr[11:4] | tagVMem_140; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_398 = 8'h8d == masterReg_Addr[11:4] | tagVMem_141; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_399 = 8'h8e == masterReg_Addr[11:4] | tagVMem_142; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_400 = 8'h8f == masterReg_Addr[11:4] | tagVMem_143; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_401 = 8'h90 == masterReg_Addr[11:4] | tagVMem_144; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_402 = 8'h91 == masterReg_Addr[11:4] | tagVMem_145; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_403 = 8'h92 == masterReg_Addr[11:4] | tagVMem_146; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_404 = 8'h93 == masterReg_Addr[11:4] | tagVMem_147; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_405 = 8'h94 == masterReg_Addr[11:4] | tagVMem_148; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_406 = 8'h95 == masterReg_Addr[11:4] | tagVMem_149; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_407 = 8'h96 == masterReg_Addr[11:4] | tagVMem_150; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_408 = 8'h97 == masterReg_Addr[11:4] | tagVMem_151; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_409 = 8'h98 == masterReg_Addr[11:4] | tagVMem_152; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_410 = 8'h99 == masterReg_Addr[11:4] | tagVMem_153; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_411 = 8'h9a == masterReg_Addr[11:4] | tagVMem_154; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_412 = 8'h9b == masterReg_Addr[11:4] | tagVMem_155; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_413 = 8'h9c == masterReg_Addr[11:4] | tagVMem_156; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_414 = 8'h9d == masterReg_Addr[11:4] | tagVMem_157; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_415 = 8'h9e == masterReg_Addr[11:4] | tagVMem_158; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_416 = 8'h9f == masterReg_Addr[11:4] | tagVMem_159; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_417 = 8'ha0 == masterReg_Addr[11:4] | tagVMem_160; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_418 = 8'ha1 == masterReg_Addr[11:4] | tagVMem_161; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_419 = 8'ha2 == masterReg_Addr[11:4] | tagVMem_162; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_420 = 8'ha3 == masterReg_Addr[11:4] | tagVMem_163; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_421 = 8'ha4 == masterReg_Addr[11:4] | tagVMem_164; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_422 = 8'ha5 == masterReg_Addr[11:4] | tagVMem_165; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_423 = 8'ha6 == masterReg_Addr[11:4] | tagVMem_166; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_424 = 8'ha7 == masterReg_Addr[11:4] | tagVMem_167; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_425 = 8'ha8 == masterReg_Addr[11:4] | tagVMem_168; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_426 = 8'ha9 == masterReg_Addr[11:4] | tagVMem_169; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_427 = 8'haa == masterReg_Addr[11:4] | tagVMem_170; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_428 = 8'hab == masterReg_Addr[11:4] | tagVMem_171; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_429 = 8'hac == masterReg_Addr[11:4] | tagVMem_172; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_430 = 8'had == masterReg_Addr[11:4] | tagVMem_173; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_431 = 8'hae == masterReg_Addr[11:4] | tagVMem_174; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_432 = 8'haf == masterReg_Addr[11:4] | tagVMem_175; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_433 = 8'hb0 == masterReg_Addr[11:4] | tagVMem_176; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_434 = 8'hb1 == masterReg_Addr[11:4] | tagVMem_177; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_435 = 8'hb2 == masterReg_Addr[11:4] | tagVMem_178; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_436 = 8'hb3 == masterReg_Addr[11:4] | tagVMem_179; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_437 = 8'hb4 == masterReg_Addr[11:4] | tagVMem_180; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_438 = 8'hb5 == masterReg_Addr[11:4] | tagVMem_181; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_439 = 8'hb6 == masterReg_Addr[11:4] | tagVMem_182; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_440 = 8'hb7 == masterReg_Addr[11:4] | tagVMem_183; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_441 = 8'hb8 == masterReg_Addr[11:4] | tagVMem_184; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_442 = 8'hb9 == masterReg_Addr[11:4] | tagVMem_185; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_443 = 8'hba == masterReg_Addr[11:4] | tagVMem_186; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_444 = 8'hbb == masterReg_Addr[11:4] | tagVMem_187; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_445 = 8'hbc == masterReg_Addr[11:4] | tagVMem_188; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_446 = 8'hbd == masterReg_Addr[11:4] | tagVMem_189; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_447 = 8'hbe == masterReg_Addr[11:4] | tagVMem_190; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_448 = 8'hbf == masterReg_Addr[11:4] | tagVMem_191; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_449 = 8'hc0 == masterReg_Addr[11:4] | tagVMem_192; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_450 = 8'hc1 == masterReg_Addr[11:4] | tagVMem_193; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_451 = 8'hc2 == masterReg_Addr[11:4] | tagVMem_194; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_452 = 8'hc3 == masterReg_Addr[11:4] | tagVMem_195; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_453 = 8'hc4 == masterReg_Addr[11:4] | tagVMem_196; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_454 = 8'hc5 == masterReg_Addr[11:4] | tagVMem_197; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_455 = 8'hc6 == masterReg_Addr[11:4] | tagVMem_198; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_456 = 8'hc7 == masterReg_Addr[11:4] | tagVMem_199; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_457 = 8'hc8 == masterReg_Addr[11:4] | tagVMem_200; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_458 = 8'hc9 == masterReg_Addr[11:4] | tagVMem_201; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_459 = 8'hca == masterReg_Addr[11:4] | tagVMem_202; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_460 = 8'hcb == masterReg_Addr[11:4] | tagVMem_203; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_461 = 8'hcc == masterReg_Addr[11:4] | tagVMem_204; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_462 = 8'hcd == masterReg_Addr[11:4] | tagVMem_205; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_463 = 8'hce == masterReg_Addr[11:4] | tagVMem_206; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_464 = 8'hcf == masterReg_Addr[11:4] | tagVMem_207; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_465 = 8'hd0 == masterReg_Addr[11:4] | tagVMem_208; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_466 = 8'hd1 == masterReg_Addr[11:4] | tagVMem_209; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_467 = 8'hd2 == masterReg_Addr[11:4] | tagVMem_210; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_468 = 8'hd3 == masterReg_Addr[11:4] | tagVMem_211; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_469 = 8'hd4 == masterReg_Addr[11:4] | tagVMem_212; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_470 = 8'hd5 == masterReg_Addr[11:4] | tagVMem_213; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_471 = 8'hd6 == masterReg_Addr[11:4] | tagVMem_214; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_472 = 8'hd7 == masterReg_Addr[11:4] | tagVMem_215; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_473 = 8'hd8 == masterReg_Addr[11:4] | tagVMem_216; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_474 = 8'hd9 == masterReg_Addr[11:4] | tagVMem_217; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_475 = 8'hda == masterReg_Addr[11:4] | tagVMem_218; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_476 = 8'hdb == masterReg_Addr[11:4] | tagVMem_219; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_477 = 8'hdc == masterReg_Addr[11:4] | tagVMem_220; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_478 = 8'hdd == masterReg_Addr[11:4] | tagVMem_221; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_479 = 8'hde == masterReg_Addr[11:4] | tagVMem_222; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_480 = 8'hdf == masterReg_Addr[11:4] | tagVMem_223; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_481 = 8'he0 == masterReg_Addr[11:4] | tagVMem_224; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_482 = 8'he1 == masterReg_Addr[11:4] | tagVMem_225; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_483 = 8'he2 == masterReg_Addr[11:4] | tagVMem_226; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_484 = 8'he3 == masterReg_Addr[11:4] | tagVMem_227; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_485 = 8'he4 == masterReg_Addr[11:4] | tagVMem_228; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_486 = 8'he5 == masterReg_Addr[11:4] | tagVMem_229; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_487 = 8'he6 == masterReg_Addr[11:4] | tagVMem_230; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_488 = 8'he7 == masterReg_Addr[11:4] | tagVMem_231; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_489 = 8'he8 == masterReg_Addr[11:4] | tagVMem_232; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_490 = 8'he9 == masterReg_Addr[11:4] | tagVMem_233; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_491 = 8'hea == masterReg_Addr[11:4] | tagVMem_234; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_492 = 8'heb == masterReg_Addr[11:4] | tagVMem_235; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_493 = 8'hec == masterReg_Addr[11:4] | tagVMem_236; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_494 = 8'hed == masterReg_Addr[11:4] | tagVMem_237; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_495 = 8'hee == masterReg_Addr[11:4] | tagVMem_238; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_496 = 8'hef == masterReg_Addr[11:4] | tagVMem_239; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_497 = 8'hf0 == masterReg_Addr[11:4] | tagVMem_240; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_498 = 8'hf1 == masterReg_Addr[11:4] | tagVMem_241; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_499 = 8'hf2 == masterReg_Addr[11:4] | tagVMem_242; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_500 = 8'hf3 == masterReg_Addr[11:4] | tagVMem_243; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_501 = 8'hf4 == masterReg_Addr[11:4] | tagVMem_244; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_502 = 8'hf5 == masterReg_Addr[11:4] | tagVMem_245; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_503 = 8'hf6 == masterReg_Addr[11:4] | tagVMem_246; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_504 = 8'hf7 == masterReg_Addr[11:4] | tagVMem_247; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_505 = 8'hf8 == masterReg_Addr[11:4] | tagVMem_248; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_506 = 8'hf9 == masterReg_Addr[11:4] | tagVMem_249; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_507 = 8'hfa == masterReg_Addr[11:4] | tagVMem_250; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_508 = 8'hfb == masterReg_Addr[11:4] | tagVMem_251; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_509 = 8'hfc == masterReg_Addr[11:4] | tagVMem_252; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_510 = 8'hfd == masterReg_Addr[11:4] | tagVMem_253; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_511 = 8'hfe == masterReg_Addr[11:4] | tagVMem_254; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire  _GEN_512 = 8'hff == masterReg_Addr[11:4] | tagVMem_255; // @[DirectMappedCache.scala 102:53 DirectMappedCache.scala 102:53 DirectMappedCache.scala 42:24]
  wire [1:0] _GEN_513 = io_slave_S_CmdAccept ? 2'h2 : 2'h1; // @[DirectMappedCache.scala 105:44 DirectMappedCache.scala 106:16 DirectMappedCache.scala 109:16]
  wire  _GEN_514 = ~tagValid & _T_28 ? _GEN_257 : tagVMem_0; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_515 = ~tagValid & _T_28 ? _GEN_258 : tagVMem_1; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_516 = ~tagValid & _T_28 ? _GEN_259 : tagVMem_2; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_517 = ~tagValid & _T_28 ? _GEN_260 : tagVMem_3; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_518 = ~tagValid & _T_28 ? _GEN_261 : tagVMem_4; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_519 = ~tagValid & _T_28 ? _GEN_262 : tagVMem_5; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_520 = ~tagValid & _T_28 ? _GEN_263 : tagVMem_6; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_521 = ~tagValid & _T_28 ? _GEN_264 : tagVMem_7; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_522 = ~tagValid & _T_28 ? _GEN_265 : tagVMem_8; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_523 = ~tagValid & _T_28 ? _GEN_266 : tagVMem_9; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_524 = ~tagValid & _T_28 ? _GEN_267 : tagVMem_10; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_525 = ~tagValid & _T_28 ? _GEN_268 : tagVMem_11; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_526 = ~tagValid & _T_28 ? _GEN_269 : tagVMem_12; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_527 = ~tagValid & _T_28 ? _GEN_270 : tagVMem_13; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_528 = ~tagValid & _T_28 ? _GEN_271 : tagVMem_14; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_529 = ~tagValid & _T_28 ? _GEN_272 : tagVMem_15; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_530 = ~tagValid & _T_28 ? _GEN_273 : tagVMem_16; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_531 = ~tagValid & _T_28 ? _GEN_274 : tagVMem_17; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_532 = ~tagValid & _T_28 ? _GEN_275 : tagVMem_18; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_533 = ~tagValid & _T_28 ? _GEN_276 : tagVMem_19; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_534 = ~tagValid & _T_28 ? _GEN_277 : tagVMem_20; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_535 = ~tagValid & _T_28 ? _GEN_278 : tagVMem_21; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_536 = ~tagValid & _T_28 ? _GEN_279 : tagVMem_22; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_537 = ~tagValid & _T_28 ? _GEN_280 : tagVMem_23; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_538 = ~tagValid & _T_28 ? _GEN_281 : tagVMem_24; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_539 = ~tagValid & _T_28 ? _GEN_282 : tagVMem_25; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_540 = ~tagValid & _T_28 ? _GEN_283 : tagVMem_26; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_541 = ~tagValid & _T_28 ? _GEN_284 : tagVMem_27; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_542 = ~tagValid & _T_28 ? _GEN_285 : tagVMem_28; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_543 = ~tagValid & _T_28 ? _GEN_286 : tagVMem_29; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_544 = ~tagValid & _T_28 ? _GEN_287 : tagVMem_30; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_545 = ~tagValid & _T_28 ? _GEN_288 : tagVMem_31; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_546 = ~tagValid & _T_28 ? _GEN_289 : tagVMem_32; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_547 = ~tagValid & _T_28 ? _GEN_290 : tagVMem_33; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_548 = ~tagValid & _T_28 ? _GEN_291 : tagVMem_34; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_549 = ~tagValid & _T_28 ? _GEN_292 : tagVMem_35; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_550 = ~tagValid & _T_28 ? _GEN_293 : tagVMem_36; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_551 = ~tagValid & _T_28 ? _GEN_294 : tagVMem_37; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_552 = ~tagValid & _T_28 ? _GEN_295 : tagVMem_38; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_553 = ~tagValid & _T_28 ? _GEN_296 : tagVMem_39; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_554 = ~tagValid & _T_28 ? _GEN_297 : tagVMem_40; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_555 = ~tagValid & _T_28 ? _GEN_298 : tagVMem_41; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_556 = ~tagValid & _T_28 ? _GEN_299 : tagVMem_42; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_557 = ~tagValid & _T_28 ? _GEN_300 : tagVMem_43; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_558 = ~tagValid & _T_28 ? _GEN_301 : tagVMem_44; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_559 = ~tagValid & _T_28 ? _GEN_302 : tagVMem_45; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_560 = ~tagValid & _T_28 ? _GEN_303 : tagVMem_46; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_561 = ~tagValid & _T_28 ? _GEN_304 : tagVMem_47; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_562 = ~tagValid & _T_28 ? _GEN_305 : tagVMem_48; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_563 = ~tagValid & _T_28 ? _GEN_306 : tagVMem_49; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_564 = ~tagValid & _T_28 ? _GEN_307 : tagVMem_50; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_565 = ~tagValid & _T_28 ? _GEN_308 : tagVMem_51; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_566 = ~tagValid & _T_28 ? _GEN_309 : tagVMem_52; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_567 = ~tagValid & _T_28 ? _GEN_310 : tagVMem_53; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_568 = ~tagValid & _T_28 ? _GEN_311 : tagVMem_54; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_569 = ~tagValid & _T_28 ? _GEN_312 : tagVMem_55; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_570 = ~tagValid & _T_28 ? _GEN_313 : tagVMem_56; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_571 = ~tagValid & _T_28 ? _GEN_314 : tagVMem_57; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_572 = ~tagValid & _T_28 ? _GEN_315 : tagVMem_58; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_573 = ~tagValid & _T_28 ? _GEN_316 : tagVMem_59; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_574 = ~tagValid & _T_28 ? _GEN_317 : tagVMem_60; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_575 = ~tagValid & _T_28 ? _GEN_318 : tagVMem_61; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_576 = ~tagValid & _T_28 ? _GEN_319 : tagVMem_62; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_577 = ~tagValid & _T_28 ? _GEN_320 : tagVMem_63; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_578 = ~tagValid & _T_28 ? _GEN_321 : tagVMem_64; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_579 = ~tagValid & _T_28 ? _GEN_322 : tagVMem_65; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_580 = ~tagValid & _T_28 ? _GEN_323 : tagVMem_66; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_581 = ~tagValid & _T_28 ? _GEN_324 : tagVMem_67; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_582 = ~tagValid & _T_28 ? _GEN_325 : tagVMem_68; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_583 = ~tagValid & _T_28 ? _GEN_326 : tagVMem_69; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_584 = ~tagValid & _T_28 ? _GEN_327 : tagVMem_70; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_585 = ~tagValid & _T_28 ? _GEN_328 : tagVMem_71; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_586 = ~tagValid & _T_28 ? _GEN_329 : tagVMem_72; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_587 = ~tagValid & _T_28 ? _GEN_330 : tagVMem_73; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_588 = ~tagValid & _T_28 ? _GEN_331 : tagVMem_74; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_589 = ~tagValid & _T_28 ? _GEN_332 : tagVMem_75; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_590 = ~tagValid & _T_28 ? _GEN_333 : tagVMem_76; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_591 = ~tagValid & _T_28 ? _GEN_334 : tagVMem_77; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_592 = ~tagValid & _T_28 ? _GEN_335 : tagVMem_78; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_593 = ~tagValid & _T_28 ? _GEN_336 : tagVMem_79; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_594 = ~tagValid & _T_28 ? _GEN_337 : tagVMem_80; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_595 = ~tagValid & _T_28 ? _GEN_338 : tagVMem_81; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_596 = ~tagValid & _T_28 ? _GEN_339 : tagVMem_82; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_597 = ~tagValid & _T_28 ? _GEN_340 : tagVMem_83; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_598 = ~tagValid & _T_28 ? _GEN_341 : tagVMem_84; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_599 = ~tagValid & _T_28 ? _GEN_342 : tagVMem_85; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_600 = ~tagValid & _T_28 ? _GEN_343 : tagVMem_86; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_601 = ~tagValid & _T_28 ? _GEN_344 : tagVMem_87; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_602 = ~tagValid & _T_28 ? _GEN_345 : tagVMem_88; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_603 = ~tagValid & _T_28 ? _GEN_346 : tagVMem_89; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_604 = ~tagValid & _T_28 ? _GEN_347 : tagVMem_90; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_605 = ~tagValid & _T_28 ? _GEN_348 : tagVMem_91; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_606 = ~tagValid & _T_28 ? _GEN_349 : tagVMem_92; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_607 = ~tagValid & _T_28 ? _GEN_350 : tagVMem_93; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_608 = ~tagValid & _T_28 ? _GEN_351 : tagVMem_94; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_609 = ~tagValid & _T_28 ? _GEN_352 : tagVMem_95; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_610 = ~tagValid & _T_28 ? _GEN_353 : tagVMem_96; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_611 = ~tagValid & _T_28 ? _GEN_354 : tagVMem_97; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_612 = ~tagValid & _T_28 ? _GEN_355 : tagVMem_98; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_613 = ~tagValid & _T_28 ? _GEN_356 : tagVMem_99; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_614 = ~tagValid & _T_28 ? _GEN_357 : tagVMem_100; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_615 = ~tagValid & _T_28 ? _GEN_358 : tagVMem_101; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_616 = ~tagValid & _T_28 ? _GEN_359 : tagVMem_102; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_617 = ~tagValid & _T_28 ? _GEN_360 : tagVMem_103; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_618 = ~tagValid & _T_28 ? _GEN_361 : tagVMem_104; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_619 = ~tagValid & _T_28 ? _GEN_362 : tagVMem_105; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_620 = ~tagValid & _T_28 ? _GEN_363 : tagVMem_106; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_621 = ~tagValid & _T_28 ? _GEN_364 : tagVMem_107; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_622 = ~tagValid & _T_28 ? _GEN_365 : tagVMem_108; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_623 = ~tagValid & _T_28 ? _GEN_366 : tagVMem_109; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_624 = ~tagValid & _T_28 ? _GEN_367 : tagVMem_110; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_625 = ~tagValid & _T_28 ? _GEN_368 : tagVMem_111; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_626 = ~tagValid & _T_28 ? _GEN_369 : tagVMem_112; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_627 = ~tagValid & _T_28 ? _GEN_370 : tagVMem_113; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_628 = ~tagValid & _T_28 ? _GEN_371 : tagVMem_114; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_629 = ~tagValid & _T_28 ? _GEN_372 : tagVMem_115; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_630 = ~tagValid & _T_28 ? _GEN_373 : tagVMem_116; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_631 = ~tagValid & _T_28 ? _GEN_374 : tagVMem_117; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_632 = ~tagValid & _T_28 ? _GEN_375 : tagVMem_118; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_633 = ~tagValid & _T_28 ? _GEN_376 : tagVMem_119; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_634 = ~tagValid & _T_28 ? _GEN_377 : tagVMem_120; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_635 = ~tagValid & _T_28 ? _GEN_378 : tagVMem_121; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_636 = ~tagValid & _T_28 ? _GEN_379 : tagVMem_122; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_637 = ~tagValid & _T_28 ? _GEN_380 : tagVMem_123; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_638 = ~tagValid & _T_28 ? _GEN_381 : tagVMem_124; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_639 = ~tagValid & _T_28 ? _GEN_382 : tagVMem_125; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_640 = ~tagValid & _T_28 ? _GEN_383 : tagVMem_126; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_641 = ~tagValid & _T_28 ? _GEN_384 : tagVMem_127; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_642 = ~tagValid & _T_28 ? _GEN_385 : tagVMem_128; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_643 = ~tagValid & _T_28 ? _GEN_386 : tagVMem_129; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_644 = ~tagValid & _T_28 ? _GEN_387 : tagVMem_130; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_645 = ~tagValid & _T_28 ? _GEN_388 : tagVMem_131; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_646 = ~tagValid & _T_28 ? _GEN_389 : tagVMem_132; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_647 = ~tagValid & _T_28 ? _GEN_390 : tagVMem_133; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_648 = ~tagValid & _T_28 ? _GEN_391 : tagVMem_134; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_649 = ~tagValid & _T_28 ? _GEN_392 : tagVMem_135; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_650 = ~tagValid & _T_28 ? _GEN_393 : tagVMem_136; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_651 = ~tagValid & _T_28 ? _GEN_394 : tagVMem_137; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_652 = ~tagValid & _T_28 ? _GEN_395 : tagVMem_138; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_653 = ~tagValid & _T_28 ? _GEN_396 : tagVMem_139; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_654 = ~tagValid & _T_28 ? _GEN_397 : tagVMem_140; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_655 = ~tagValid & _T_28 ? _GEN_398 : tagVMem_141; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_656 = ~tagValid & _T_28 ? _GEN_399 : tagVMem_142; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_657 = ~tagValid & _T_28 ? _GEN_400 : tagVMem_143; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_658 = ~tagValid & _T_28 ? _GEN_401 : tagVMem_144; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_659 = ~tagValid & _T_28 ? _GEN_402 : tagVMem_145; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_660 = ~tagValid & _T_28 ? _GEN_403 : tagVMem_146; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_661 = ~tagValid & _T_28 ? _GEN_404 : tagVMem_147; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_662 = ~tagValid & _T_28 ? _GEN_405 : tagVMem_148; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_663 = ~tagValid & _T_28 ? _GEN_406 : tagVMem_149; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_664 = ~tagValid & _T_28 ? _GEN_407 : tagVMem_150; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_665 = ~tagValid & _T_28 ? _GEN_408 : tagVMem_151; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_666 = ~tagValid & _T_28 ? _GEN_409 : tagVMem_152; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_667 = ~tagValid & _T_28 ? _GEN_410 : tagVMem_153; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_668 = ~tagValid & _T_28 ? _GEN_411 : tagVMem_154; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_669 = ~tagValid & _T_28 ? _GEN_412 : tagVMem_155; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_670 = ~tagValid & _T_28 ? _GEN_413 : tagVMem_156; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_671 = ~tagValid & _T_28 ? _GEN_414 : tagVMem_157; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_672 = ~tagValid & _T_28 ? _GEN_415 : tagVMem_158; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_673 = ~tagValid & _T_28 ? _GEN_416 : tagVMem_159; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_674 = ~tagValid & _T_28 ? _GEN_417 : tagVMem_160; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_675 = ~tagValid & _T_28 ? _GEN_418 : tagVMem_161; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_676 = ~tagValid & _T_28 ? _GEN_419 : tagVMem_162; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_677 = ~tagValid & _T_28 ? _GEN_420 : tagVMem_163; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_678 = ~tagValid & _T_28 ? _GEN_421 : tagVMem_164; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_679 = ~tagValid & _T_28 ? _GEN_422 : tagVMem_165; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_680 = ~tagValid & _T_28 ? _GEN_423 : tagVMem_166; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_681 = ~tagValid & _T_28 ? _GEN_424 : tagVMem_167; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_682 = ~tagValid & _T_28 ? _GEN_425 : tagVMem_168; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_683 = ~tagValid & _T_28 ? _GEN_426 : tagVMem_169; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_684 = ~tagValid & _T_28 ? _GEN_427 : tagVMem_170; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_685 = ~tagValid & _T_28 ? _GEN_428 : tagVMem_171; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_686 = ~tagValid & _T_28 ? _GEN_429 : tagVMem_172; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_687 = ~tagValid & _T_28 ? _GEN_430 : tagVMem_173; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_688 = ~tagValid & _T_28 ? _GEN_431 : tagVMem_174; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_689 = ~tagValid & _T_28 ? _GEN_432 : tagVMem_175; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_690 = ~tagValid & _T_28 ? _GEN_433 : tagVMem_176; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_691 = ~tagValid & _T_28 ? _GEN_434 : tagVMem_177; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_692 = ~tagValid & _T_28 ? _GEN_435 : tagVMem_178; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_693 = ~tagValid & _T_28 ? _GEN_436 : tagVMem_179; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_694 = ~tagValid & _T_28 ? _GEN_437 : tagVMem_180; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_695 = ~tagValid & _T_28 ? _GEN_438 : tagVMem_181; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_696 = ~tagValid & _T_28 ? _GEN_439 : tagVMem_182; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_697 = ~tagValid & _T_28 ? _GEN_440 : tagVMem_183; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_698 = ~tagValid & _T_28 ? _GEN_441 : tagVMem_184; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_699 = ~tagValid & _T_28 ? _GEN_442 : tagVMem_185; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_700 = ~tagValid & _T_28 ? _GEN_443 : tagVMem_186; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_701 = ~tagValid & _T_28 ? _GEN_444 : tagVMem_187; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_702 = ~tagValid & _T_28 ? _GEN_445 : tagVMem_188; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_703 = ~tagValid & _T_28 ? _GEN_446 : tagVMem_189; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_704 = ~tagValid & _T_28 ? _GEN_447 : tagVMem_190; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_705 = ~tagValid & _T_28 ? _GEN_448 : tagVMem_191; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_706 = ~tagValid & _T_28 ? _GEN_449 : tagVMem_192; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_707 = ~tagValid & _T_28 ? _GEN_450 : tagVMem_193; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_708 = ~tagValid & _T_28 ? _GEN_451 : tagVMem_194; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_709 = ~tagValid & _T_28 ? _GEN_452 : tagVMem_195; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_710 = ~tagValid & _T_28 ? _GEN_453 : tagVMem_196; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_711 = ~tagValid & _T_28 ? _GEN_454 : tagVMem_197; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_712 = ~tagValid & _T_28 ? _GEN_455 : tagVMem_198; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_713 = ~tagValid & _T_28 ? _GEN_456 : tagVMem_199; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_714 = ~tagValid & _T_28 ? _GEN_457 : tagVMem_200; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_715 = ~tagValid & _T_28 ? _GEN_458 : tagVMem_201; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_716 = ~tagValid & _T_28 ? _GEN_459 : tagVMem_202; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_717 = ~tagValid & _T_28 ? _GEN_460 : tagVMem_203; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_718 = ~tagValid & _T_28 ? _GEN_461 : tagVMem_204; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_719 = ~tagValid & _T_28 ? _GEN_462 : tagVMem_205; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_720 = ~tagValid & _T_28 ? _GEN_463 : tagVMem_206; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_721 = ~tagValid & _T_28 ? _GEN_464 : tagVMem_207; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_722 = ~tagValid & _T_28 ? _GEN_465 : tagVMem_208; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_723 = ~tagValid & _T_28 ? _GEN_466 : tagVMem_209; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_724 = ~tagValid & _T_28 ? _GEN_467 : tagVMem_210; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_725 = ~tagValid & _T_28 ? _GEN_468 : tagVMem_211; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_726 = ~tagValid & _T_28 ? _GEN_469 : tagVMem_212; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_727 = ~tagValid & _T_28 ? _GEN_470 : tagVMem_213; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_728 = ~tagValid & _T_28 ? _GEN_471 : tagVMem_214; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_729 = ~tagValid & _T_28 ? _GEN_472 : tagVMem_215; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_730 = ~tagValid & _T_28 ? _GEN_473 : tagVMem_216; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_731 = ~tagValid & _T_28 ? _GEN_474 : tagVMem_217; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_732 = ~tagValid & _T_28 ? _GEN_475 : tagVMem_218; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_733 = ~tagValid & _T_28 ? _GEN_476 : tagVMem_219; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_734 = ~tagValid & _T_28 ? _GEN_477 : tagVMem_220; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_735 = ~tagValid & _T_28 ? _GEN_478 : tagVMem_221; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_736 = ~tagValid & _T_28 ? _GEN_479 : tagVMem_222; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_737 = ~tagValid & _T_28 ? _GEN_480 : tagVMem_223; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_738 = ~tagValid & _T_28 ? _GEN_481 : tagVMem_224; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_739 = ~tagValid & _T_28 ? _GEN_482 : tagVMem_225; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_740 = ~tagValid & _T_28 ? _GEN_483 : tagVMem_226; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_741 = ~tagValid & _T_28 ? _GEN_484 : tagVMem_227; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_742 = ~tagValid & _T_28 ? _GEN_485 : tagVMem_228; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_743 = ~tagValid & _T_28 ? _GEN_486 : tagVMem_229; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_744 = ~tagValid & _T_28 ? _GEN_487 : tagVMem_230; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_745 = ~tagValid & _T_28 ? _GEN_488 : tagVMem_231; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_746 = ~tagValid & _T_28 ? _GEN_489 : tagVMem_232; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_747 = ~tagValid & _T_28 ? _GEN_490 : tagVMem_233; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_748 = ~tagValid & _T_28 ? _GEN_491 : tagVMem_234; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_749 = ~tagValid & _T_28 ? _GEN_492 : tagVMem_235; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_750 = ~tagValid & _T_28 ? _GEN_493 : tagVMem_236; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_751 = ~tagValid & _T_28 ? _GEN_494 : tagVMem_237; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_752 = ~tagValid & _T_28 ? _GEN_495 : tagVMem_238; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_753 = ~tagValid & _T_28 ? _GEN_496 : tagVMem_239; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_754 = ~tagValid & _T_28 ? _GEN_497 : tagVMem_240; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_755 = ~tagValid & _T_28 ? _GEN_498 : tagVMem_241; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_756 = ~tagValid & _T_28 ? _GEN_499 : tagVMem_242; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_757 = ~tagValid & _T_28 ? _GEN_500 : tagVMem_243; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_758 = ~tagValid & _T_28 ? _GEN_501 : tagVMem_244; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_759 = ~tagValid & _T_28 ? _GEN_502 : tagVMem_245; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_760 = ~tagValid & _T_28 ? _GEN_503 : tagVMem_246; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_761 = ~tagValid & _T_28 ? _GEN_504 : tagVMem_247; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_762 = ~tagValid & _T_28 ? _GEN_505 : tagVMem_248; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_763 = ~tagValid & _T_28 ? _GEN_506 : tagVMem_249; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_764 = ~tagValid & _T_28 ? _GEN_507 : tagVMem_250; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_765 = ~tagValid & _T_28 ? _GEN_508 : tagVMem_251; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_766 = ~tagValid & _T_28 ? _GEN_509 : tagVMem_252; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_767 = ~tagValid & _T_28 ? _GEN_510 : tagVMem_253; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_768 = ~tagValid & _T_28 ? _GEN_511 : tagVMem_254; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire  _GEN_769 = ~tagValid & _T_28 ? _GEN_512 : tagVMem_255; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 42:24]
  wire [2:0] _GEN_771 = ~tagValid & _T_28 ? 3'h2 : 3'h0; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 104:20 DirectMappedCache.scala 86:18]
  wire [1:0] _GEN_772 = ~tagValid & _T_28 ? _GEN_513 : stateReg; // @[DirectMappedCache.scala 101:50 DirectMappedCache.scala 77:21]
  wire [1:0] _GEN_777 = stateReg == 2'h1 ? _GEN_513 : _GEN_772; // @[DirectMappedCache.scala 119:27]
  wire [9:0] _T_48 = {masterReg_Addr[11:4],burstCntReg}; // @[Cat.scala 30:58]
  wire  _T_49 = io_slave_S_Resp != 2'h0; // @[DirectMappedCache.scala 133:26]
  wire [1:0] _GEN_781 = burstCntReg == 2'h3 ? 2'h3 : _GEN_777; // @[DirectMappedCache.scala 139:48 DirectMappedCache.scala 140:18]
  wire [1:0] _lo_T_1 = burstCntReg + 2'h1; // @[DirectMappedCache.scala 142:34]
  wire  _GEN_788 = 8'h0 == masterReg_Addr[11:4] ? 1'h0 : _GEN_514; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_789 = 8'h1 == masterReg_Addr[11:4] ? 1'h0 : _GEN_515; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_790 = 8'h2 == masterReg_Addr[11:4] ? 1'h0 : _GEN_516; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_791 = 8'h3 == masterReg_Addr[11:4] ? 1'h0 : _GEN_517; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_792 = 8'h4 == masterReg_Addr[11:4] ? 1'h0 : _GEN_518; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_793 = 8'h5 == masterReg_Addr[11:4] ? 1'h0 : _GEN_519; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_794 = 8'h6 == masterReg_Addr[11:4] ? 1'h0 : _GEN_520; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_795 = 8'h7 == masterReg_Addr[11:4] ? 1'h0 : _GEN_521; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_796 = 8'h8 == masterReg_Addr[11:4] ? 1'h0 : _GEN_522; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_797 = 8'h9 == masterReg_Addr[11:4] ? 1'h0 : _GEN_523; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_798 = 8'ha == masterReg_Addr[11:4] ? 1'h0 : _GEN_524; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_799 = 8'hb == masterReg_Addr[11:4] ? 1'h0 : _GEN_525; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_800 = 8'hc == masterReg_Addr[11:4] ? 1'h0 : _GEN_526; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_801 = 8'hd == masterReg_Addr[11:4] ? 1'h0 : _GEN_527; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_802 = 8'he == masterReg_Addr[11:4] ? 1'h0 : _GEN_528; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_803 = 8'hf == masterReg_Addr[11:4] ? 1'h0 : _GEN_529; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_804 = 8'h10 == masterReg_Addr[11:4] ? 1'h0 : _GEN_530; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_805 = 8'h11 == masterReg_Addr[11:4] ? 1'h0 : _GEN_531; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_806 = 8'h12 == masterReg_Addr[11:4] ? 1'h0 : _GEN_532; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_807 = 8'h13 == masterReg_Addr[11:4] ? 1'h0 : _GEN_533; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_808 = 8'h14 == masterReg_Addr[11:4] ? 1'h0 : _GEN_534; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_809 = 8'h15 == masterReg_Addr[11:4] ? 1'h0 : _GEN_535; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_810 = 8'h16 == masterReg_Addr[11:4] ? 1'h0 : _GEN_536; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_811 = 8'h17 == masterReg_Addr[11:4] ? 1'h0 : _GEN_537; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_812 = 8'h18 == masterReg_Addr[11:4] ? 1'h0 : _GEN_538; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_813 = 8'h19 == masterReg_Addr[11:4] ? 1'h0 : _GEN_539; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_814 = 8'h1a == masterReg_Addr[11:4] ? 1'h0 : _GEN_540; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_815 = 8'h1b == masterReg_Addr[11:4] ? 1'h0 : _GEN_541; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_816 = 8'h1c == masterReg_Addr[11:4] ? 1'h0 : _GEN_542; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_817 = 8'h1d == masterReg_Addr[11:4] ? 1'h0 : _GEN_543; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_818 = 8'h1e == masterReg_Addr[11:4] ? 1'h0 : _GEN_544; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_819 = 8'h1f == masterReg_Addr[11:4] ? 1'h0 : _GEN_545; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_820 = 8'h20 == masterReg_Addr[11:4] ? 1'h0 : _GEN_546; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_821 = 8'h21 == masterReg_Addr[11:4] ? 1'h0 : _GEN_547; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_822 = 8'h22 == masterReg_Addr[11:4] ? 1'h0 : _GEN_548; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_823 = 8'h23 == masterReg_Addr[11:4] ? 1'h0 : _GEN_549; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_824 = 8'h24 == masterReg_Addr[11:4] ? 1'h0 : _GEN_550; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_825 = 8'h25 == masterReg_Addr[11:4] ? 1'h0 : _GEN_551; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_826 = 8'h26 == masterReg_Addr[11:4] ? 1'h0 : _GEN_552; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_827 = 8'h27 == masterReg_Addr[11:4] ? 1'h0 : _GEN_553; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_828 = 8'h28 == masterReg_Addr[11:4] ? 1'h0 : _GEN_554; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_829 = 8'h29 == masterReg_Addr[11:4] ? 1'h0 : _GEN_555; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_830 = 8'h2a == masterReg_Addr[11:4] ? 1'h0 : _GEN_556; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_831 = 8'h2b == masterReg_Addr[11:4] ? 1'h0 : _GEN_557; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_832 = 8'h2c == masterReg_Addr[11:4] ? 1'h0 : _GEN_558; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_833 = 8'h2d == masterReg_Addr[11:4] ? 1'h0 : _GEN_559; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_834 = 8'h2e == masterReg_Addr[11:4] ? 1'h0 : _GEN_560; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_835 = 8'h2f == masterReg_Addr[11:4] ? 1'h0 : _GEN_561; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_836 = 8'h30 == masterReg_Addr[11:4] ? 1'h0 : _GEN_562; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_837 = 8'h31 == masterReg_Addr[11:4] ? 1'h0 : _GEN_563; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_838 = 8'h32 == masterReg_Addr[11:4] ? 1'h0 : _GEN_564; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_839 = 8'h33 == masterReg_Addr[11:4] ? 1'h0 : _GEN_565; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_840 = 8'h34 == masterReg_Addr[11:4] ? 1'h0 : _GEN_566; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_841 = 8'h35 == masterReg_Addr[11:4] ? 1'h0 : _GEN_567; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_842 = 8'h36 == masterReg_Addr[11:4] ? 1'h0 : _GEN_568; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_843 = 8'h37 == masterReg_Addr[11:4] ? 1'h0 : _GEN_569; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_844 = 8'h38 == masterReg_Addr[11:4] ? 1'h0 : _GEN_570; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_845 = 8'h39 == masterReg_Addr[11:4] ? 1'h0 : _GEN_571; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_846 = 8'h3a == masterReg_Addr[11:4] ? 1'h0 : _GEN_572; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_847 = 8'h3b == masterReg_Addr[11:4] ? 1'h0 : _GEN_573; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_848 = 8'h3c == masterReg_Addr[11:4] ? 1'h0 : _GEN_574; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_849 = 8'h3d == masterReg_Addr[11:4] ? 1'h0 : _GEN_575; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_850 = 8'h3e == masterReg_Addr[11:4] ? 1'h0 : _GEN_576; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_851 = 8'h3f == masterReg_Addr[11:4] ? 1'h0 : _GEN_577; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_852 = 8'h40 == masterReg_Addr[11:4] ? 1'h0 : _GEN_578; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_853 = 8'h41 == masterReg_Addr[11:4] ? 1'h0 : _GEN_579; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_854 = 8'h42 == masterReg_Addr[11:4] ? 1'h0 : _GEN_580; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_855 = 8'h43 == masterReg_Addr[11:4] ? 1'h0 : _GEN_581; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_856 = 8'h44 == masterReg_Addr[11:4] ? 1'h0 : _GEN_582; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_857 = 8'h45 == masterReg_Addr[11:4] ? 1'h0 : _GEN_583; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_858 = 8'h46 == masterReg_Addr[11:4] ? 1'h0 : _GEN_584; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_859 = 8'h47 == masterReg_Addr[11:4] ? 1'h0 : _GEN_585; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_860 = 8'h48 == masterReg_Addr[11:4] ? 1'h0 : _GEN_586; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_861 = 8'h49 == masterReg_Addr[11:4] ? 1'h0 : _GEN_587; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_862 = 8'h4a == masterReg_Addr[11:4] ? 1'h0 : _GEN_588; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_863 = 8'h4b == masterReg_Addr[11:4] ? 1'h0 : _GEN_589; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_864 = 8'h4c == masterReg_Addr[11:4] ? 1'h0 : _GEN_590; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_865 = 8'h4d == masterReg_Addr[11:4] ? 1'h0 : _GEN_591; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_866 = 8'h4e == masterReg_Addr[11:4] ? 1'h0 : _GEN_592; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_867 = 8'h4f == masterReg_Addr[11:4] ? 1'h0 : _GEN_593; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_868 = 8'h50 == masterReg_Addr[11:4] ? 1'h0 : _GEN_594; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_869 = 8'h51 == masterReg_Addr[11:4] ? 1'h0 : _GEN_595; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_870 = 8'h52 == masterReg_Addr[11:4] ? 1'h0 : _GEN_596; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_871 = 8'h53 == masterReg_Addr[11:4] ? 1'h0 : _GEN_597; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_872 = 8'h54 == masterReg_Addr[11:4] ? 1'h0 : _GEN_598; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_873 = 8'h55 == masterReg_Addr[11:4] ? 1'h0 : _GEN_599; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_874 = 8'h56 == masterReg_Addr[11:4] ? 1'h0 : _GEN_600; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_875 = 8'h57 == masterReg_Addr[11:4] ? 1'h0 : _GEN_601; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_876 = 8'h58 == masterReg_Addr[11:4] ? 1'h0 : _GEN_602; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_877 = 8'h59 == masterReg_Addr[11:4] ? 1'h0 : _GEN_603; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_878 = 8'h5a == masterReg_Addr[11:4] ? 1'h0 : _GEN_604; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_879 = 8'h5b == masterReg_Addr[11:4] ? 1'h0 : _GEN_605; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_880 = 8'h5c == masterReg_Addr[11:4] ? 1'h0 : _GEN_606; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_881 = 8'h5d == masterReg_Addr[11:4] ? 1'h0 : _GEN_607; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_882 = 8'h5e == masterReg_Addr[11:4] ? 1'h0 : _GEN_608; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_883 = 8'h5f == masterReg_Addr[11:4] ? 1'h0 : _GEN_609; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_884 = 8'h60 == masterReg_Addr[11:4] ? 1'h0 : _GEN_610; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_885 = 8'h61 == masterReg_Addr[11:4] ? 1'h0 : _GEN_611; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_886 = 8'h62 == masterReg_Addr[11:4] ? 1'h0 : _GEN_612; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_887 = 8'h63 == masterReg_Addr[11:4] ? 1'h0 : _GEN_613; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_888 = 8'h64 == masterReg_Addr[11:4] ? 1'h0 : _GEN_614; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_889 = 8'h65 == masterReg_Addr[11:4] ? 1'h0 : _GEN_615; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_890 = 8'h66 == masterReg_Addr[11:4] ? 1'h0 : _GEN_616; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_891 = 8'h67 == masterReg_Addr[11:4] ? 1'h0 : _GEN_617; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_892 = 8'h68 == masterReg_Addr[11:4] ? 1'h0 : _GEN_618; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_893 = 8'h69 == masterReg_Addr[11:4] ? 1'h0 : _GEN_619; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_894 = 8'h6a == masterReg_Addr[11:4] ? 1'h0 : _GEN_620; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_895 = 8'h6b == masterReg_Addr[11:4] ? 1'h0 : _GEN_621; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_896 = 8'h6c == masterReg_Addr[11:4] ? 1'h0 : _GEN_622; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_897 = 8'h6d == masterReg_Addr[11:4] ? 1'h0 : _GEN_623; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_898 = 8'h6e == masterReg_Addr[11:4] ? 1'h0 : _GEN_624; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_899 = 8'h6f == masterReg_Addr[11:4] ? 1'h0 : _GEN_625; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_900 = 8'h70 == masterReg_Addr[11:4] ? 1'h0 : _GEN_626; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_901 = 8'h71 == masterReg_Addr[11:4] ? 1'h0 : _GEN_627; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_902 = 8'h72 == masterReg_Addr[11:4] ? 1'h0 : _GEN_628; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_903 = 8'h73 == masterReg_Addr[11:4] ? 1'h0 : _GEN_629; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_904 = 8'h74 == masterReg_Addr[11:4] ? 1'h0 : _GEN_630; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_905 = 8'h75 == masterReg_Addr[11:4] ? 1'h0 : _GEN_631; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_906 = 8'h76 == masterReg_Addr[11:4] ? 1'h0 : _GEN_632; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_907 = 8'h77 == masterReg_Addr[11:4] ? 1'h0 : _GEN_633; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_908 = 8'h78 == masterReg_Addr[11:4] ? 1'h0 : _GEN_634; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_909 = 8'h79 == masterReg_Addr[11:4] ? 1'h0 : _GEN_635; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_910 = 8'h7a == masterReg_Addr[11:4] ? 1'h0 : _GEN_636; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_911 = 8'h7b == masterReg_Addr[11:4] ? 1'h0 : _GEN_637; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_912 = 8'h7c == masterReg_Addr[11:4] ? 1'h0 : _GEN_638; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_913 = 8'h7d == masterReg_Addr[11:4] ? 1'h0 : _GEN_639; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_914 = 8'h7e == masterReg_Addr[11:4] ? 1'h0 : _GEN_640; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_915 = 8'h7f == masterReg_Addr[11:4] ? 1'h0 : _GEN_641; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_916 = 8'h80 == masterReg_Addr[11:4] ? 1'h0 : _GEN_642; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_917 = 8'h81 == masterReg_Addr[11:4] ? 1'h0 : _GEN_643; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_918 = 8'h82 == masterReg_Addr[11:4] ? 1'h0 : _GEN_644; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_919 = 8'h83 == masterReg_Addr[11:4] ? 1'h0 : _GEN_645; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_920 = 8'h84 == masterReg_Addr[11:4] ? 1'h0 : _GEN_646; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_921 = 8'h85 == masterReg_Addr[11:4] ? 1'h0 : _GEN_647; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_922 = 8'h86 == masterReg_Addr[11:4] ? 1'h0 : _GEN_648; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_923 = 8'h87 == masterReg_Addr[11:4] ? 1'h0 : _GEN_649; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_924 = 8'h88 == masterReg_Addr[11:4] ? 1'h0 : _GEN_650; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_925 = 8'h89 == masterReg_Addr[11:4] ? 1'h0 : _GEN_651; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_926 = 8'h8a == masterReg_Addr[11:4] ? 1'h0 : _GEN_652; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_927 = 8'h8b == masterReg_Addr[11:4] ? 1'h0 : _GEN_653; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_928 = 8'h8c == masterReg_Addr[11:4] ? 1'h0 : _GEN_654; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_929 = 8'h8d == masterReg_Addr[11:4] ? 1'h0 : _GEN_655; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_930 = 8'h8e == masterReg_Addr[11:4] ? 1'h0 : _GEN_656; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_931 = 8'h8f == masterReg_Addr[11:4] ? 1'h0 : _GEN_657; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_932 = 8'h90 == masterReg_Addr[11:4] ? 1'h0 : _GEN_658; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_933 = 8'h91 == masterReg_Addr[11:4] ? 1'h0 : _GEN_659; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_934 = 8'h92 == masterReg_Addr[11:4] ? 1'h0 : _GEN_660; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_935 = 8'h93 == masterReg_Addr[11:4] ? 1'h0 : _GEN_661; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_936 = 8'h94 == masterReg_Addr[11:4] ? 1'h0 : _GEN_662; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_937 = 8'h95 == masterReg_Addr[11:4] ? 1'h0 : _GEN_663; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_938 = 8'h96 == masterReg_Addr[11:4] ? 1'h0 : _GEN_664; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_939 = 8'h97 == masterReg_Addr[11:4] ? 1'h0 : _GEN_665; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_940 = 8'h98 == masterReg_Addr[11:4] ? 1'h0 : _GEN_666; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_941 = 8'h99 == masterReg_Addr[11:4] ? 1'h0 : _GEN_667; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_942 = 8'h9a == masterReg_Addr[11:4] ? 1'h0 : _GEN_668; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_943 = 8'h9b == masterReg_Addr[11:4] ? 1'h0 : _GEN_669; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_944 = 8'h9c == masterReg_Addr[11:4] ? 1'h0 : _GEN_670; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_945 = 8'h9d == masterReg_Addr[11:4] ? 1'h0 : _GEN_671; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_946 = 8'h9e == masterReg_Addr[11:4] ? 1'h0 : _GEN_672; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_947 = 8'h9f == masterReg_Addr[11:4] ? 1'h0 : _GEN_673; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_948 = 8'ha0 == masterReg_Addr[11:4] ? 1'h0 : _GEN_674; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_949 = 8'ha1 == masterReg_Addr[11:4] ? 1'h0 : _GEN_675; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_950 = 8'ha2 == masterReg_Addr[11:4] ? 1'h0 : _GEN_676; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_951 = 8'ha3 == masterReg_Addr[11:4] ? 1'h0 : _GEN_677; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_952 = 8'ha4 == masterReg_Addr[11:4] ? 1'h0 : _GEN_678; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_953 = 8'ha5 == masterReg_Addr[11:4] ? 1'h0 : _GEN_679; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_954 = 8'ha6 == masterReg_Addr[11:4] ? 1'h0 : _GEN_680; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_955 = 8'ha7 == masterReg_Addr[11:4] ? 1'h0 : _GEN_681; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_956 = 8'ha8 == masterReg_Addr[11:4] ? 1'h0 : _GEN_682; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_957 = 8'ha9 == masterReg_Addr[11:4] ? 1'h0 : _GEN_683; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_958 = 8'haa == masterReg_Addr[11:4] ? 1'h0 : _GEN_684; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_959 = 8'hab == masterReg_Addr[11:4] ? 1'h0 : _GEN_685; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_960 = 8'hac == masterReg_Addr[11:4] ? 1'h0 : _GEN_686; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_961 = 8'had == masterReg_Addr[11:4] ? 1'h0 : _GEN_687; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_962 = 8'hae == masterReg_Addr[11:4] ? 1'h0 : _GEN_688; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_963 = 8'haf == masterReg_Addr[11:4] ? 1'h0 : _GEN_689; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_964 = 8'hb0 == masterReg_Addr[11:4] ? 1'h0 : _GEN_690; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_965 = 8'hb1 == masterReg_Addr[11:4] ? 1'h0 : _GEN_691; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_966 = 8'hb2 == masterReg_Addr[11:4] ? 1'h0 : _GEN_692; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_967 = 8'hb3 == masterReg_Addr[11:4] ? 1'h0 : _GEN_693; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_968 = 8'hb4 == masterReg_Addr[11:4] ? 1'h0 : _GEN_694; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_969 = 8'hb5 == masterReg_Addr[11:4] ? 1'h0 : _GEN_695; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_970 = 8'hb6 == masterReg_Addr[11:4] ? 1'h0 : _GEN_696; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_971 = 8'hb7 == masterReg_Addr[11:4] ? 1'h0 : _GEN_697; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_972 = 8'hb8 == masterReg_Addr[11:4] ? 1'h0 : _GEN_698; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_973 = 8'hb9 == masterReg_Addr[11:4] ? 1'h0 : _GEN_699; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_974 = 8'hba == masterReg_Addr[11:4] ? 1'h0 : _GEN_700; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_975 = 8'hbb == masterReg_Addr[11:4] ? 1'h0 : _GEN_701; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_976 = 8'hbc == masterReg_Addr[11:4] ? 1'h0 : _GEN_702; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_977 = 8'hbd == masterReg_Addr[11:4] ? 1'h0 : _GEN_703; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_978 = 8'hbe == masterReg_Addr[11:4] ? 1'h0 : _GEN_704; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_979 = 8'hbf == masterReg_Addr[11:4] ? 1'h0 : _GEN_705; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_980 = 8'hc0 == masterReg_Addr[11:4] ? 1'h0 : _GEN_706; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_981 = 8'hc1 == masterReg_Addr[11:4] ? 1'h0 : _GEN_707; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_982 = 8'hc2 == masterReg_Addr[11:4] ? 1'h0 : _GEN_708; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_983 = 8'hc3 == masterReg_Addr[11:4] ? 1'h0 : _GEN_709; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_984 = 8'hc4 == masterReg_Addr[11:4] ? 1'h0 : _GEN_710; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_985 = 8'hc5 == masterReg_Addr[11:4] ? 1'h0 : _GEN_711; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_986 = 8'hc6 == masterReg_Addr[11:4] ? 1'h0 : _GEN_712; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_987 = 8'hc7 == masterReg_Addr[11:4] ? 1'h0 : _GEN_713; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_988 = 8'hc8 == masterReg_Addr[11:4] ? 1'h0 : _GEN_714; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_989 = 8'hc9 == masterReg_Addr[11:4] ? 1'h0 : _GEN_715; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_990 = 8'hca == masterReg_Addr[11:4] ? 1'h0 : _GEN_716; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_991 = 8'hcb == masterReg_Addr[11:4] ? 1'h0 : _GEN_717; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_992 = 8'hcc == masterReg_Addr[11:4] ? 1'h0 : _GEN_718; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_993 = 8'hcd == masterReg_Addr[11:4] ? 1'h0 : _GEN_719; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_994 = 8'hce == masterReg_Addr[11:4] ? 1'h0 : _GEN_720; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_995 = 8'hcf == masterReg_Addr[11:4] ? 1'h0 : _GEN_721; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_996 = 8'hd0 == masterReg_Addr[11:4] ? 1'h0 : _GEN_722; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_997 = 8'hd1 == masterReg_Addr[11:4] ? 1'h0 : _GEN_723; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_998 = 8'hd2 == masterReg_Addr[11:4] ? 1'h0 : _GEN_724; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_999 = 8'hd3 == masterReg_Addr[11:4] ? 1'h0 : _GEN_725; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1000 = 8'hd4 == masterReg_Addr[11:4] ? 1'h0 : _GEN_726; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1001 = 8'hd5 == masterReg_Addr[11:4] ? 1'h0 : _GEN_727; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1002 = 8'hd6 == masterReg_Addr[11:4] ? 1'h0 : _GEN_728; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1003 = 8'hd7 == masterReg_Addr[11:4] ? 1'h0 : _GEN_729; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1004 = 8'hd8 == masterReg_Addr[11:4] ? 1'h0 : _GEN_730; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1005 = 8'hd9 == masterReg_Addr[11:4] ? 1'h0 : _GEN_731; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1006 = 8'hda == masterReg_Addr[11:4] ? 1'h0 : _GEN_732; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1007 = 8'hdb == masterReg_Addr[11:4] ? 1'h0 : _GEN_733; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1008 = 8'hdc == masterReg_Addr[11:4] ? 1'h0 : _GEN_734; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1009 = 8'hdd == masterReg_Addr[11:4] ? 1'h0 : _GEN_735; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1010 = 8'hde == masterReg_Addr[11:4] ? 1'h0 : _GEN_736; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1011 = 8'hdf == masterReg_Addr[11:4] ? 1'h0 : _GEN_737; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1012 = 8'he0 == masterReg_Addr[11:4] ? 1'h0 : _GEN_738; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1013 = 8'he1 == masterReg_Addr[11:4] ? 1'h0 : _GEN_739; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1014 = 8'he2 == masterReg_Addr[11:4] ? 1'h0 : _GEN_740; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1015 = 8'he3 == masterReg_Addr[11:4] ? 1'h0 : _GEN_741; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1016 = 8'he4 == masterReg_Addr[11:4] ? 1'h0 : _GEN_742; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1017 = 8'he5 == masterReg_Addr[11:4] ? 1'h0 : _GEN_743; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1018 = 8'he6 == masterReg_Addr[11:4] ? 1'h0 : _GEN_744; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1019 = 8'he7 == masterReg_Addr[11:4] ? 1'h0 : _GEN_745; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1020 = 8'he8 == masterReg_Addr[11:4] ? 1'h0 : _GEN_746; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1021 = 8'he9 == masterReg_Addr[11:4] ? 1'h0 : _GEN_747; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1022 = 8'hea == masterReg_Addr[11:4] ? 1'h0 : _GEN_748; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1023 = 8'heb == masterReg_Addr[11:4] ? 1'h0 : _GEN_749; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1024 = 8'hec == masterReg_Addr[11:4] ? 1'h0 : _GEN_750; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1025 = 8'hed == masterReg_Addr[11:4] ? 1'h0 : _GEN_751; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1026 = 8'hee == masterReg_Addr[11:4] ? 1'h0 : _GEN_752; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1027 = 8'hef == masterReg_Addr[11:4] ? 1'h0 : _GEN_753; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1028 = 8'hf0 == masterReg_Addr[11:4] ? 1'h0 : _GEN_754; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1029 = 8'hf1 == masterReg_Addr[11:4] ? 1'h0 : _GEN_755; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1030 = 8'hf2 == masterReg_Addr[11:4] ? 1'h0 : _GEN_756; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1031 = 8'hf3 == masterReg_Addr[11:4] ? 1'h0 : _GEN_757; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1032 = 8'hf4 == masterReg_Addr[11:4] ? 1'h0 : _GEN_758; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1033 = 8'hf5 == masterReg_Addr[11:4] ? 1'h0 : _GEN_759; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1034 = 8'hf6 == masterReg_Addr[11:4] ? 1'h0 : _GEN_760; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1035 = 8'hf7 == masterReg_Addr[11:4] ? 1'h0 : _GEN_761; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1036 = 8'hf8 == masterReg_Addr[11:4] ? 1'h0 : _GEN_762; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1037 = 8'hf9 == masterReg_Addr[11:4] ? 1'h0 : _GEN_763; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1038 = 8'hfa == masterReg_Addr[11:4] ? 1'h0 : _GEN_764; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1039 = 8'hfb == masterReg_Addr[11:4] ? 1'h0 : _GEN_765; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1040 = 8'hfc == masterReg_Addr[11:4] ? 1'h0 : _GEN_766; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1041 = 8'hfd == masterReg_Addr[11:4] ? 1'h0 : _GEN_767; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1042 = 8'hfe == masterReg_Addr[11:4] ? 1'h0 : _GEN_768; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  wire  _GEN_1043 = 8'hff == masterReg_Addr[11:4] ? 1'h0 : _GEN_769; // @[DirectMappedCache.scala 145:55 DirectMappedCache.scala 145:55]
  MemBlock_4 tagMem ( // @[MemBlock.scala 15:11]
    .clock(tagMem_clock),
    .io_rdAddr(tagMem_io_rdAddr),
    .io_rdData(tagMem_io_rdData),
    .io_wrAddr(tagMem_io_wrAddr),
    .io_wrEna(tagMem_io_wrEna),
    .io_wrData(tagMem_io_wrData)
  );
  MemBlock_5 MemBlock ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_clock),
    .io_rdAddr(MemBlock_io_rdAddr),
    .io_rdData(MemBlock_io_rdData),
    .io_wrAddr(MemBlock_io_wrAddr),
    .io_wrEna(MemBlock_io_wrEna),
    .io_wrData(MemBlock_io_wrData)
  );
  MemBlock_5 MemBlock_1 ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_1_clock),
    .io_rdAddr(MemBlock_1_io_rdAddr),
    .io_rdData(MemBlock_1_io_rdData),
    .io_wrAddr(MemBlock_1_io_wrAddr),
    .io_wrEna(MemBlock_1_io_wrEna),
    .io_wrData(MemBlock_1_io_wrData)
  );
  MemBlock_5 MemBlock_2 ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_2_clock),
    .io_rdAddr(MemBlock_2_io_rdAddr),
    .io_rdData(MemBlock_2_io_rdData),
    .io_wrAddr(MemBlock_2_io_wrAddr),
    .io_wrEna(MemBlock_2_io_wrEna),
    .io_wrData(MemBlock_2_io_wrData)
  );
  MemBlock_5 MemBlock_3 ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_3_clock),
    .io_rdAddr(MemBlock_3_io_rdAddr),
    .io_rdData(MemBlock_3_io_rdData),
    .io_wrAddr(MemBlock_3_io_wrAddr),
    .io_wrEna(MemBlock_3_io_wrEna),
    .io_wrData(MemBlock_3_io_wrData)
  );
  assign io_master_S_Resp = stateReg == 2'h3 ? slaveReg_Resp : _T_30; // @[DirectMappedCache.scala 150:30 DirectMappedCache.scala 151:17 DirectMappedCache.scala 72:20]
  assign io_master_S_Data = stateReg == 2'h3 ? slaveReg_Data : rdData; // @[DirectMappedCache.scala 150:30 DirectMappedCache.scala 151:17 DirectMappedCache.scala 71:20]
  assign io_slave_M_Cmd = stateReg == 2'h1 ? 3'h2 : _GEN_771; // @[DirectMappedCache.scala 119:27 DirectMappedCache.scala 120:20]
  assign io_slave_M_Addr = {hi,4'h0}; // @[Cat.scala 30:58]
  assign tagMem_clock = clock;
  assign tagMem_io_rdAddr = io_master_M_Addr[11:4]; // @[DirectMappedCache.scala 48:39]
  assign tagMem_io_wrAddr = masterReg_Addr[11:4]; // @[DirectMappedCache.scala 115:31]
  assign tagMem_io_wrEna = _T_34 & _T_28; // @[DirectMappedCache.scala 114:27]
  assign tagMem_io_wrData = masterReg_Addr[31:12]; // @[DirectMappedCache.scala 116:31]
  assign MemBlock_clock = clock;
  assign MemBlock_io_rdAddr = io_master_M_Addr[11:2]; // @[DirectMappedCache.scala 68:42]
  assign MemBlock_io_wrAddr = wrAddrReg; // @[MemBlock.scala 34:12]
  assign MemBlock_io_wrEna = fillReg | tagValid & stmsk[0]; // @[DirectMappedCache.scala 63:24]
  assign MemBlock_io_wrData = wrDataReg[7:0]; // @[DirectMappedCache.scala 64:25]
  assign MemBlock_1_clock = clock;
  assign MemBlock_1_io_rdAddr = io_master_M_Addr[11:2]; // @[DirectMappedCache.scala 68:42]
  assign MemBlock_1_io_wrAddr = wrAddrReg; // @[MemBlock.scala 34:12]
  assign MemBlock_1_io_wrEna = fillReg | tagValid & stmsk[1]; // @[DirectMappedCache.scala 63:24]
  assign MemBlock_1_io_wrData = wrDataReg[15:8]; // @[DirectMappedCache.scala 64:25]
  assign MemBlock_2_clock = clock;
  assign MemBlock_2_io_rdAddr = io_master_M_Addr[11:2]; // @[DirectMappedCache.scala 68:42]
  assign MemBlock_2_io_wrAddr = wrAddrReg; // @[MemBlock.scala 34:12]
  assign MemBlock_2_io_wrEna = fillReg | tagValid & stmsk[2]; // @[DirectMappedCache.scala 63:24]
  assign MemBlock_2_io_wrData = wrDataReg[23:16]; // @[DirectMappedCache.scala 64:25]
  assign MemBlock_3_clock = clock;
  assign MemBlock_3_io_rdAddr = io_master_M_Addr[11:2]; // @[DirectMappedCache.scala 68:42]
  assign MemBlock_3_io_wrAddr = wrAddrReg; // @[MemBlock.scala 34:12]
  assign MemBlock_3_io_wrEna = fillReg | tagValid & stmsk[3]; // @[DirectMappedCache.scala 63:24]
  assign MemBlock_3_io_wrData = wrDataReg[31:24]; // @[DirectMappedCache.scala 64:25]
  always @(posedge clock) begin
    masterReg_Cmd <= io_master_M_Cmd; // @[DirectMappedCache.scala 38:13]
    if (!(stateReg == 2'h2)) begin // @[DirectMappedCache.scala 130:27]
      if (!(stateReg == 2'h1)) begin // @[DirectMappedCache.scala 119:27]
        if (!(~tagValid & _T_28)) begin // @[DirectMappedCache.scala 101:50]
          masterReg_Addr <= io_master_M_Addr; // @[DirectMappedCache.scala 38:13]
        end
      end
    end
    masterReg_ByteEn <= io_master_M_ByteEn; // @[DirectMappedCache.scala 38:13]
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_0 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_0 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_0 <= _GEN_788;
      end else begin
        tagVMem_0 <= _GEN_514;
      end
    end else begin
      tagVMem_0 <= _GEN_514;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_1 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_1 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_1 <= _GEN_789;
      end else begin
        tagVMem_1 <= _GEN_515;
      end
    end else begin
      tagVMem_1 <= _GEN_515;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_2 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_2 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_2 <= _GEN_790;
      end else begin
        tagVMem_2 <= _GEN_516;
      end
    end else begin
      tagVMem_2 <= _GEN_516;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_3 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_3 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_3 <= _GEN_791;
      end else begin
        tagVMem_3 <= _GEN_517;
      end
    end else begin
      tagVMem_3 <= _GEN_517;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_4 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_4 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_4 <= _GEN_792;
      end else begin
        tagVMem_4 <= _GEN_518;
      end
    end else begin
      tagVMem_4 <= _GEN_518;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_5 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_5 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_5 <= _GEN_793;
      end else begin
        tagVMem_5 <= _GEN_519;
      end
    end else begin
      tagVMem_5 <= _GEN_519;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_6 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_6 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_6 <= _GEN_794;
      end else begin
        tagVMem_6 <= _GEN_520;
      end
    end else begin
      tagVMem_6 <= _GEN_520;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_7 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_7 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_7 <= _GEN_795;
      end else begin
        tagVMem_7 <= _GEN_521;
      end
    end else begin
      tagVMem_7 <= _GEN_521;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_8 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_8 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_8 <= _GEN_796;
      end else begin
        tagVMem_8 <= _GEN_522;
      end
    end else begin
      tagVMem_8 <= _GEN_522;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_9 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_9 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_9 <= _GEN_797;
      end else begin
        tagVMem_9 <= _GEN_523;
      end
    end else begin
      tagVMem_9 <= _GEN_523;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_10 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_10 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_10 <= _GEN_798;
      end else begin
        tagVMem_10 <= _GEN_524;
      end
    end else begin
      tagVMem_10 <= _GEN_524;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_11 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_11 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_11 <= _GEN_799;
      end else begin
        tagVMem_11 <= _GEN_525;
      end
    end else begin
      tagVMem_11 <= _GEN_525;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_12 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_12 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_12 <= _GEN_800;
      end else begin
        tagVMem_12 <= _GEN_526;
      end
    end else begin
      tagVMem_12 <= _GEN_526;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_13 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_13 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_13 <= _GEN_801;
      end else begin
        tagVMem_13 <= _GEN_527;
      end
    end else begin
      tagVMem_13 <= _GEN_527;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_14 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_14 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_14 <= _GEN_802;
      end else begin
        tagVMem_14 <= _GEN_528;
      end
    end else begin
      tagVMem_14 <= _GEN_528;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_15 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_15 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_15 <= _GEN_803;
      end else begin
        tagVMem_15 <= _GEN_529;
      end
    end else begin
      tagVMem_15 <= _GEN_529;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_16 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_16 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_16 <= _GEN_804;
      end else begin
        tagVMem_16 <= _GEN_530;
      end
    end else begin
      tagVMem_16 <= _GEN_530;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_17 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_17 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_17 <= _GEN_805;
      end else begin
        tagVMem_17 <= _GEN_531;
      end
    end else begin
      tagVMem_17 <= _GEN_531;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_18 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_18 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_18 <= _GEN_806;
      end else begin
        tagVMem_18 <= _GEN_532;
      end
    end else begin
      tagVMem_18 <= _GEN_532;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_19 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_19 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_19 <= _GEN_807;
      end else begin
        tagVMem_19 <= _GEN_533;
      end
    end else begin
      tagVMem_19 <= _GEN_533;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_20 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_20 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_20 <= _GEN_808;
      end else begin
        tagVMem_20 <= _GEN_534;
      end
    end else begin
      tagVMem_20 <= _GEN_534;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_21 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_21 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_21 <= _GEN_809;
      end else begin
        tagVMem_21 <= _GEN_535;
      end
    end else begin
      tagVMem_21 <= _GEN_535;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_22 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_22 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_22 <= _GEN_810;
      end else begin
        tagVMem_22 <= _GEN_536;
      end
    end else begin
      tagVMem_22 <= _GEN_536;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_23 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_23 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_23 <= _GEN_811;
      end else begin
        tagVMem_23 <= _GEN_537;
      end
    end else begin
      tagVMem_23 <= _GEN_537;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_24 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_24 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_24 <= _GEN_812;
      end else begin
        tagVMem_24 <= _GEN_538;
      end
    end else begin
      tagVMem_24 <= _GEN_538;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_25 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_25 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_25 <= _GEN_813;
      end else begin
        tagVMem_25 <= _GEN_539;
      end
    end else begin
      tagVMem_25 <= _GEN_539;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_26 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_26 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_26 <= _GEN_814;
      end else begin
        tagVMem_26 <= _GEN_540;
      end
    end else begin
      tagVMem_26 <= _GEN_540;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_27 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_27 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_27 <= _GEN_815;
      end else begin
        tagVMem_27 <= _GEN_541;
      end
    end else begin
      tagVMem_27 <= _GEN_541;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_28 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_28 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_28 <= _GEN_816;
      end else begin
        tagVMem_28 <= _GEN_542;
      end
    end else begin
      tagVMem_28 <= _GEN_542;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_29 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_29 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_29 <= _GEN_817;
      end else begin
        tagVMem_29 <= _GEN_543;
      end
    end else begin
      tagVMem_29 <= _GEN_543;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_30 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_30 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_30 <= _GEN_818;
      end else begin
        tagVMem_30 <= _GEN_544;
      end
    end else begin
      tagVMem_30 <= _GEN_544;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_31 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_31 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_31 <= _GEN_819;
      end else begin
        tagVMem_31 <= _GEN_545;
      end
    end else begin
      tagVMem_31 <= _GEN_545;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_32 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_32 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_32 <= _GEN_820;
      end else begin
        tagVMem_32 <= _GEN_546;
      end
    end else begin
      tagVMem_32 <= _GEN_546;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_33 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_33 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_33 <= _GEN_821;
      end else begin
        tagVMem_33 <= _GEN_547;
      end
    end else begin
      tagVMem_33 <= _GEN_547;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_34 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_34 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_34 <= _GEN_822;
      end else begin
        tagVMem_34 <= _GEN_548;
      end
    end else begin
      tagVMem_34 <= _GEN_548;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_35 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_35 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_35 <= _GEN_823;
      end else begin
        tagVMem_35 <= _GEN_549;
      end
    end else begin
      tagVMem_35 <= _GEN_549;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_36 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_36 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_36 <= _GEN_824;
      end else begin
        tagVMem_36 <= _GEN_550;
      end
    end else begin
      tagVMem_36 <= _GEN_550;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_37 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_37 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_37 <= _GEN_825;
      end else begin
        tagVMem_37 <= _GEN_551;
      end
    end else begin
      tagVMem_37 <= _GEN_551;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_38 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_38 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_38 <= _GEN_826;
      end else begin
        tagVMem_38 <= _GEN_552;
      end
    end else begin
      tagVMem_38 <= _GEN_552;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_39 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_39 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_39 <= _GEN_827;
      end else begin
        tagVMem_39 <= _GEN_553;
      end
    end else begin
      tagVMem_39 <= _GEN_553;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_40 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_40 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_40 <= _GEN_828;
      end else begin
        tagVMem_40 <= _GEN_554;
      end
    end else begin
      tagVMem_40 <= _GEN_554;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_41 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_41 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_41 <= _GEN_829;
      end else begin
        tagVMem_41 <= _GEN_555;
      end
    end else begin
      tagVMem_41 <= _GEN_555;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_42 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_42 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_42 <= _GEN_830;
      end else begin
        tagVMem_42 <= _GEN_556;
      end
    end else begin
      tagVMem_42 <= _GEN_556;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_43 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_43 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_43 <= _GEN_831;
      end else begin
        tagVMem_43 <= _GEN_557;
      end
    end else begin
      tagVMem_43 <= _GEN_557;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_44 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_44 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_44 <= _GEN_832;
      end else begin
        tagVMem_44 <= _GEN_558;
      end
    end else begin
      tagVMem_44 <= _GEN_558;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_45 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_45 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_45 <= _GEN_833;
      end else begin
        tagVMem_45 <= _GEN_559;
      end
    end else begin
      tagVMem_45 <= _GEN_559;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_46 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_46 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_46 <= _GEN_834;
      end else begin
        tagVMem_46 <= _GEN_560;
      end
    end else begin
      tagVMem_46 <= _GEN_560;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_47 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_47 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_47 <= _GEN_835;
      end else begin
        tagVMem_47 <= _GEN_561;
      end
    end else begin
      tagVMem_47 <= _GEN_561;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_48 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_48 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_48 <= _GEN_836;
      end else begin
        tagVMem_48 <= _GEN_562;
      end
    end else begin
      tagVMem_48 <= _GEN_562;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_49 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_49 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_49 <= _GEN_837;
      end else begin
        tagVMem_49 <= _GEN_563;
      end
    end else begin
      tagVMem_49 <= _GEN_563;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_50 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_50 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_50 <= _GEN_838;
      end else begin
        tagVMem_50 <= _GEN_564;
      end
    end else begin
      tagVMem_50 <= _GEN_564;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_51 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_51 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_51 <= _GEN_839;
      end else begin
        tagVMem_51 <= _GEN_565;
      end
    end else begin
      tagVMem_51 <= _GEN_565;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_52 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_52 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_52 <= _GEN_840;
      end else begin
        tagVMem_52 <= _GEN_566;
      end
    end else begin
      tagVMem_52 <= _GEN_566;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_53 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_53 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_53 <= _GEN_841;
      end else begin
        tagVMem_53 <= _GEN_567;
      end
    end else begin
      tagVMem_53 <= _GEN_567;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_54 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_54 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_54 <= _GEN_842;
      end else begin
        tagVMem_54 <= _GEN_568;
      end
    end else begin
      tagVMem_54 <= _GEN_568;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_55 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_55 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_55 <= _GEN_843;
      end else begin
        tagVMem_55 <= _GEN_569;
      end
    end else begin
      tagVMem_55 <= _GEN_569;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_56 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_56 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_56 <= _GEN_844;
      end else begin
        tagVMem_56 <= _GEN_570;
      end
    end else begin
      tagVMem_56 <= _GEN_570;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_57 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_57 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_57 <= _GEN_845;
      end else begin
        tagVMem_57 <= _GEN_571;
      end
    end else begin
      tagVMem_57 <= _GEN_571;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_58 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_58 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_58 <= _GEN_846;
      end else begin
        tagVMem_58 <= _GEN_572;
      end
    end else begin
      tagVMem_58 <= _GEN_572;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_59 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_59 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_59 <= _GEN_847;
      end else begin
        tagVMem_59 <= _GEN_573;
      end
    end else begin
      tagVMem_59 <= _GEN_573;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_60 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_60 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_60 <= _GEN_848;
      end else begin
        tagVMem_60 <= _GEN_574;
      end
    end else begin
      tagVMem_60 <= _GEN_574;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_61 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_61 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_61 <= _GEN_849;
      end else begin
        tagVMem_61 <= _GEN_575;
      end
    end else begin
      tagVMem_61 <= _GEN_575;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_62 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_62 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_62 <= _GEN_850;
      end else begin
        tagVMem_62 <= _GEN_576;
      end
    end else begin
      tagVMem_62 <= _GEN_576;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_63 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_63 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_63 <= _GEN_851;
      end else begin
        tagVMem_63 <= _GEN_577;
      end
    end else begin
      tagVMem_63 <= _GEN_577;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_64 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_64 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_64 <= _GEN_852;
      end else begin
        tagVMem_64 <= _GEN_578;
      end
    end else begin
      tagVMem_64 <= _GEN_578;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_65 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_65 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_65 <= _GEN_853;
      end else begin
        tagVMem_65 <= _GEN_579;
      end
    end else begin
      tagVMem_65 <= _GEN_579;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_66 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_66 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_66 <= _GEN_854;
      end else begin
        tagVMem_66 <= _GEN_580;
      end
    end else begin
      tagVMem_66 <= _GEN_580;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_67 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_67 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_67 <= _GEN_855;
      end else begin
        tagVMem_67 <= _GEN_581;
      end
    end else begin
      tagVMem_67 <= _GEN_581;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_68 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_68 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_68 <= _GEN_856;
      end else begin
        tagVMem_68 <= _GEN_582;
      end
    end else begin
      tagVMem_68 <= _GEN_582;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_69 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_69 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_69 <= _GEN_857;
      end else begin
        tagVMem_69 <= _GEN_583;
      end
    end else begin
      tagVMem_69 <= _GEN_583;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_70 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_70 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_70 <= _GEN_858;
      end else begin
        tagVMem_70 <= _GEN_584;
      end
    end else begin
      tagVMem_70 <= _GEN_584;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_71 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_71 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_71 <= _GEN_859;
      end else begin
        tagVMem_71 <= _GEN_585;
      end
    end else begin
      tagVMem_71 <= _GEN_585;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_72 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_72 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_72 <= _GEN_860;
      end else begin
        tagVMem_72 <= _GEN_586;
      end
    end else begin
      tagVMem_72 <= _GEN_586;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_73 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_73 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_73 <= _GEN_861;
      end else begin
        tagVMem_73 <= _GEN_587;
      end
    end else begin
      tagVMem_73 <= _GEN_587;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_74 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_74 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_74 <= _GEN_862;
      end else begin
        tagVMem_74 <= _GEN_588;
      end
    end else begin
      tagVMem_74 <= _GEN_588;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_75 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_75 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_75 <= _GEN_863;
      end else begin
        tagVMem_75 <= _GEN_589;
      end
    end else begin
      tagVMem_75 <= _GEN_589;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_76 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_76 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_76 <= _GEN_864;
      end else begin
        tagVMem_76 <= _GEN_590;
      end
    end else begin
      tagVMem_76 <= _GEN_590;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_77 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_77 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_77 <= _GEN_865;
      end else begin
        tagVMem_77 <= _GEN_591;
      end
    end else begin
      tagVMem_77 <= _GEN_591;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_78 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_78 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_78 <= _GEN_866;
      end else begin
        tagVMem_78 <= _GEN_592;
      end
    end else begin
      tagVMem_78 <= _GEN_592;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_79 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_79 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_79 <= _GEN_867;
      end else begin
        tagVMem_79 <= _GEN_593;
      end
    end else begin
      tagVMem_79 <= _GEN_593;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_80 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_80 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_80 <= _GEN_868;
      end else begin
        tagVMem_80 <= _GEN_594;
      end
    end else begin
      tagVMem_80 <= _GEN_594;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_81 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_81 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_81 <= _GEN_869;
      end else begin
        tagVMem_81 <= _GEN_595;
      end
    end else begin
      tagVMem_81 <= _GEN_595;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_82 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_82 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_82 <= _GEN_870;
      end else begin
        tagVMem_82 <= _GEN_596;
      end
    end else begin
      tagVMem_82 <= _GEN_596;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_83 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_83 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_83 <= _GEN_871;
      end else begin
        tagVMem_83 <= _GEN_597;
      end
    end else begin
      tagVMem_83 <= _GEN_597;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_84 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_84 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_84 <= _GEN_872;
      end else begin
        tagVMem_84 <= _GEN_598;
      end
    end else begin
      tagVMem_84 <= _GEN_598;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_85 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_85 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_85 <= _GEN_873;
      end else begin
        tagVMem_85 <= _GEN_599;
      end
    end else begin
      tagVMem_85 <= _GEN_599;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_86 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_86 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_86 <= _GEN_874;
      end else begin
        tagVMem_86 <= _GEN_600;
      end
    end else begin
      tagVMem_86 <= _GEN_600;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_87 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_87 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_87 <= _GEN_875;
      end else begin
        tagVMem_87 <= _GEN_601;
      end
    end else begin
      tagVMem_87 <= _GEN_601;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_88 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_88 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_88 <= _GEN_876;
      end else begin
        tagVMem_88 <= _GEN_602;
      end
    end else begin
      tagVMem_88 <= _GEN_602;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_89 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_89 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_89 <= _GEN_877;
      end else begin
        tagVMem_89 <= _GEN_603;
      end
    end else begin
      tagVMem_89 <= _GEN_603;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_90 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_90 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_90 <= _GEN_878;
      end else begin
        tagVMem_90 <= _GEN_604;
      end
    end else begin
      tagVMem_90 <= _GEN_604;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_91 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_91 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_91 <= _GEN_879;
      end else begin
        tagVMem_91 <= _GEN_605;
      end
    end else begin
      tagVMem_91 <= _GEN_605;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_92 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_92 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_92 <= _GEN_880;
      end else begin
        tagVMem_92 <= _GEN_606;
      end
    end else begin
      tagVMem_92 <= _GEN_606;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_93 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_93 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_93 <= _GEN_881;
      end else begin
        tagVMem_93 <= _GEN_607;
      end
    end else begin
      tagVMem_93 <= _GEN_607;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_94 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_94 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_94 <= _GEN_882;
      end else begin
        tagVMem_94 <= _GEN_608;
      end
    end else begin
      tagVMem_94 <= _GEN_608;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_95 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_95 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_95 <= _GEN_883;
      end else begin
        tagVMem_95 <= _GEN_609;
      end
    end else begin
      tagVMem_95 <= _GEN_609;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_96 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_96 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_96 <= _GEN_884;
      end else begin
        tagVMem_96 <= _GEN_610;
      end
    end else begin
      tagVMem_96 <= _GEN_610;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_97 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_97 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_97 <= _GEN_885;
      end else begin
        tagVMem_97 <= _GEN_611;
      end
    end else begin
      tagVMem_97 <= _GEN_611;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_98 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_98 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_98 <= _GEN_886;
      end else begin
        tagVMem_98 <= _GEN_612;
      end
    end else begin
      tagVMem_98 <= _GEN_612;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_99 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_99 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_99 <= _GEN_887;
      end else begin
        tagVMem_99 <= _GEN_613;
      end
    end else begin
      tagVMem_99 <= _GEN_613;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_100 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_100 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_100 <= _GEN_888;
      end else begin
        tagVMem_100 <= _GEN_614;
      end
    end else begin
      tagVMem_100 <= _GEN_614;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_101 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_101 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_101 <= _GEN_889;
      end else begin
        tagVMem_101 <= _GEN_615;
      end
    end else begin
      tagVMem_101 <= _GEN_615;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_102 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_102 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_102 <= _GEN_890;
      end else begin
        tagVMem_102 <= _GEN_616;
      end
    end else begin
      tagVMem_102 <= _GEN_616;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_103 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_103 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_103 <= _GEN_891;
      end else begin
        tagVMem_103 <= _GEN_617;
      end
    end else begin
      tagVMem_103 <= _GEN_617;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_104 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_104 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_104 <= _GEN_892;
      end else begin
        tagVMem_104 <= _GEN_618;
      end
    end else begin
      tagVMem_104 <= _GEN_618;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_105 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_105 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_105 <= _GEN_893;
      end else begin
        tagVMem_105 <= _GEN_619;
      end
    end else begin
      tagVMem_105 <= _GEN_619;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_106 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_106 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_106 <= _GEN_894;
      end else begin
        tagVMem_106 <= _GEN_620;
      end
    end else begin
      tagVMem_106 <= _GEN_620;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_107 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_107 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_107 <= _GEN_895;
      end else begin
        tagVMem_107 <= _GEN_621;
      end
    end else begin
      tagVMem_107 <= _GEN_621;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_108 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_108 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_108 <= _GEN_896;
      end else begin
        tagVMem_108 <= _GEN_622;
      end
    end else begin
      tagVMem_108 <= _GEN_622;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_109 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_109 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_109 <= _GEN_897;
      end else begin
        tagVMem_109 <= _GEN_623;
      end
    end else begin
      tagVMem_109 <= _GEN_623;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_110 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_110 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_110 <= _GEN_898;
      end else begin
        tagVMem_110 <= _GEN_624;
      end
    end else begin
      tagVMem_110 <= _GEN_624;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_111 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_111 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_111 <= _GEN_899;
      end else begin
        tagVMem_111 <= _GEN_625;
      end
    end else begin
      tagVMem_111 <= _GEN_625;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_112 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_112 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_112 <= _GEN_900;
      end else begin
        tagVMem_112 <= _GEN_626;
      end
    end else begin
      tagVMem_112 <= _GEN_626;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_113 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_113 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_113 <= _GEN_901;
      end else begin
        tagVMem_113 <= _GEN_627;
      end
    end else begin
      tagVMem_113 <= _GEN_627;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_114 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_114 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_114 <= _GEN_902;
      end else begin
        tagVMem_114 <= _GEN_628;
      end
    end else begin
      tagVMem_114 <= _GEN_628;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_115 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_115 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_115 <= _GEN_903;
      end else begin
        tagVMem_115 <= _GEN_629;
      end
    end else begin
      tagVMem_115 <= _GEN_629;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_116 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_116 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_116 <= _GEN_904;
      end else begin
        tagVMem_116 <= _GEN_630;
      end
    end else begin
      tagVMem_116 <= _GEN_630;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_117 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_117 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_117 <= _GEN_905;
      end else begin
        tagVMem_117 <= _GEN_631;
      end
    end else begin
      tagVMem_117 <= _GEN_631;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_118 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_118 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_118 <= _GEN_906;
      end else begin
        tagVMem_118 <= _GEN_632;
      end
    end else begin
      tagVMem_118 <= _GEN_632;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_119 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_119 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_119 <= _GEN_907;
      end else begin
        tagVMem_119 <= _GEN_633;
      end
    end else begin
      tagVMem_119 <= _GEN_633;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_120 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_120 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_120 <= _GEN_908;
      end else begin
        tagVMem_120 <= _GEN_634;
      end
    end else begin
      tagVMem_120 <= _GEN_634;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_121 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_121 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_121 <= _GEN_909;
      end else begin
        tagVMem_121 <= _GEN_635;
      end
    end else begin
      tagVMem_121 <= _GEN_635;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_122 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_122 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_122 <= _GEN_910;
      end else begin
        tagVMem_122 <= _GEN_636;
      end
    end else begin
      tagVMem_122 <= _GEN_636;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_123 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_123 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_123 <= _GEN_911;
      end else begin
        tagVMem_123 <= _GEN_637;
      end
    end else begin
      tagVMem_123 <= _GEN_637;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_124 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_124 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_124 <= _GEN_912;
      end else begin
        tagVMem_124 <= _GEN_638;
      end
    end else begin
      tagVMem_124 <= _GEN_638;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_125 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_125 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_125 <= _GEN_913;
      end else begin
        tagVMem_125 <= _GEN_639;
      end
    end else begin
      tagVMem_125 <= _GEN_639;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_126 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_126 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_126 <= _GEN_914;
      end else begin
        tagVMem_126 <= _GEN_640;
      end
    end else begin
      tagVMem_126 <= _GEN_640;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_127 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_127 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_127 <= _GEN_915;
      end else begin
        tagVMem_127 <= _GEN_641;
      end
    end else begin
      tagVMem_127 <= _GEN_641;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_128 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_128 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_128 <= _GEN_916;
      end else begin
        tagVMem_128 <= _GEN_642;
      end
    end else begin
      tagVMem_128 <= _GEN_642;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_129 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_129 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_129 <= _GEN_917;
      end else begin
        tagVMem_129 <= _GEN_643;
      end
    end else begin
      tagVMem_129 <= _GEN_643;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_130 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_130 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_130 <= _GEN_918;
      end else begin
        tagVMem_130 <= _GEN_644;
      end
    end else begin
      tagVMem_130 <= _GEN_644;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_131 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_131 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_131 <= _GEN_919;
      end else begin
        tagVMem_131 <= _GEN_645;
      end
    end else begin
      tagVMem_131 <= _GEN_645;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_132 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_132 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_132 <= _GEN_920;
      end else begin
        tagVMem_132 <= _GEN_646;
      end
    end else begin
      tagVMem_132 <= _GEN_646;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_133 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_133 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_133 <= _GEN_921;
      end else begin
        tagVMem_133 <= _GEN_647;
      end
    end else begin
      tagVMem_133 <= _GEN_647;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_134 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_134 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_134 <= _GEN_922;
      end else begin
        tagVMem_134 <= _GEN_648;
      end
    end else begin
      tagVMem_134 <= _GEN_648;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_135 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_135 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_135 <= _GEN_923;
      end else begin
        tagVMem_135 <= _GEN_649;
      end
    end else begin
      tagVMem_135 <= _GEN_649;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_136 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_136 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_136 <= _GEN_924;
      end else begin
        tagVMem_136 <= _GEN_650;
      end
    end else begin
      tagVMem_136 <= _GEN_650;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_137 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_137 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_137 <= _GEN_925;
      end else begin
        tagVMem_137 <= _GEN_651;
      end
    end else begin
      tagVMem_137 <= _GEN_651;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_138 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_138 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_138 <= _GEN_926;
      end else begin
        tagVMem_138 <= _GEN_652;
      end
    end else begin
      tagVMem_138 <= _GEN_652;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_139 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_139 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_139 <= _GEN_927;
      end else begin
        tagVMem_139 <= _GEN_653;
      end
    end else begin
      tagVMem_139 <= _GEN_653;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_140 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_140 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_140 <= _GEN_928;
      end else begin
        tagVMem_140 <= _GEN_654;
      end
    end else begin
      tagVMem_140 <= _GEN_654;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_141 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_141 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_141 <= _GEN_929;
      end else begin
        tagVMem_141 <= _GEN_655;
      end
    end else begin
      tagVMem_141 <= _GEN_655;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_142 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_142 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_142 <= _GEN_930;
      end else begin
        tagVMem_142 <= _GEN_656;
      end
    end else begin
      tagVMem_142 <= _GEN_656;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_143 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_143 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_143 <= _GEN_931;
      end else begin
        tagVMem_143 <= _GEN_657;
      end
    end else begin
      tagVMem_143 <= _GEN_657;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_144 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_144 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_144 <= _GEN_932;
      end else begin
        tagVMem_144 <= _GEN_658;
      end
    end else begin
      tagVMem_144 <= _GEN_658;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_145 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_145 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_145 <= _GEN_933;
      end else begin
        tagVMem_145 <= _GEN_659;
      end
    end else begin
      tagVMem_145 <= _GEN_659;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_146 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_146 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_146 <= _GEN_934;
      end else begin
        tagVMem_146 <= _GEN_660;
      end
    end else begin
      tagVMem_146 <= _GEN_660;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_147 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_147 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_147 <= _GEN_935;
      end else begin
        tagVMem_147 <= _GEN_661;
      end
    end else begin
      tagVMem_147 <= _GEN_661;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_148 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_148 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_148 <= _GEN_936;
      end else begin
        tagVMem_148 <= _GEN_662;
      end
    end else begin
      tagVMem_148 <= _GEN_662;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_149 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_149 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_149 <= _GEN_937;
      end else begin
        tagVMem_149 <= _GEN_663;
      end
    end else begin
      tagVMem_149 <= _GEN_663;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_150 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_150 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_150 <= _GEN_938;
      end else begin
        tagVMem_150 <= _GEN_664;
      end
    end else begin
      tagVMem_150 <= _GEN_664;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_151 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_151 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_151 <= _GEN_939;
      end else begin
        tagVMem_151 <= _GEN_665;
      end
    end else begin
      tagVMem_151 <= _GEN_665;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_152 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_152 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_152 <= _GEN_940;
      end else begin
        tagVMem_152 <= _GEN_666;
      end
    end else begin
      tagVMem_152 <= _GEN_666;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_153 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_153 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_153 <= _GEN_941;
      end else begin
        tagVMem_153 <= _GEN_667;
      end
    end else begin
      tagVMem_153 <= _GEN_667;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_154 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_154 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_154 <= _GEN_942;
      end else begin
        tagVMem_154 <= _GEN_668;
      end
    end else begin
      tagVMem_154 <= _GEN_668;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_155 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_155 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_155 <= _GEN_943;
      end else begin
        tagVMem_155 <= _GEN_669;
      end
    end else begin
      tagVMem_155 <= _GEN_669;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_156 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_156 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_156 <= _GEN_944;
      end else begin
        tagVMem_156 <= _GEN_670;
      end
    end else begin
      tagVMem_156 <= _GEN_670;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_157 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_157 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_157 <= _GEN_945;
      end else begin
        tagVMem_157 <= _GEN_671;
      end
    end else begin
      tagVMem_157 <= _GEN_671;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_158 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_158 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_158 <= _GEN_946;
      end else begin
        tagVMem_158 <= _GEN_672;
      end
    end else begin
      tagVMem_158 <= _GEN_672;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_159 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_159 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_159 <= _GEN_947;
      end else begin
        tagVMem_159 <= _GEN_673;
      end
    end else begin
      tagVMem_159 <= _GEN_673;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_160 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_160 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_160 <= _GEN_948;
      end else begin
        tagVMem_160 <= _GEN_674;
      end
    end else begin
      tagVMem_160 <= _GEN_674;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_161 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_161 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_161 <= _GEN_949;
      end else begin
        tagVMem_161 <= _GEN_675;
      end
    end else begin
      tagVMem_161 <= _GEN_675;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_162 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_162 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_162 <= _GEN_950;
      end else begin
        tagVMem_162 <= _GEN_676;
      end
    end else begin
      tagVMem_162 <= _GEN_676;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_163 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_163 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_163 <= _GEN_951;
      end else begin
        tagVMem_163 <= _GEN_677;
      end
    end else begin
      tagVMem_163 <= _GEN_677;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_164 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_164 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_164 <= _GEN_952;
      end else begin
        tagVMem_164 <= _GEN_678;
      end
    end else begin
      tagVMem_164 <= _GEN_678;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_165 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_165 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_165 <= _GEN_953;
      end else begin
        tagVMem_165 <= _GEN_679;
      end
    end else begin
      tagVMem_165 <= _GEN_679;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_166 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_166 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_166 <= _GEN_954;
      end else begin
        tagVMem_166 <= _GEN_680;
      end
    end else begin
      tagVMem_166 <= _GEN_680;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_167 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_167 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_167 <= _GEN_955;
      end else begin
        tagVMem_167 <= _GEN_681;
      end
    end else begin
      tagVMem_167 <= _GEN_681;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_168 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_168 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_168 <= _GEN_956;
      end else begin
        tagVMem_168 <= _GEN_682;
      end
    end else begin
      tagVMem_168 <= _GEN_682;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_169 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_169 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_169 <= _GEN_957;
      end else begin
        tagVMem_169 <= _GEN_683;
      end
    end else begin
      tagVMem_169 <= _GEN_683;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_170 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_170 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_170 <= _GEN_958;
      end else begin
        tagVMem_170 <= _GEN_684;
      end
    end else begin
      tagVMem_170 <= _GEN_684;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_171 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_171 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_171 <= _GEN_959;
      end else begin
        tagVMem_171 <= _GEN_685;
      end
    end else begin
      tagVMem_171 <= _GEN_685;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_172 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_172 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_172 <= _GEN_960;
      end else begin
        tagVMem_172 <= _GEN_686;
      end
    end else begin
      tagVMem_172 <= _GEN_686;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_173 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_173 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_173 <= _GEN_961;
      end else begin
        tagVMem_173 <= _GEN_687;
      end
    end else begin
      tagVMem_173 <= _GEN_687;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_174 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_174 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_174 <= _GEN_962;
      end else begin
        tagVMem_174 <= _GEN_688;
      end
    end else begin
      tagVMem_174 <= _GEN_688;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_175 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_175 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_175 <= _GEN_963;
      end else begin
        tagVMem_175 <= _GEN_689;
      end
    end else begin
      tagVMem_175 <= _GEN_689;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_176 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_176 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_176 <= _GEN_964;
      end else begin
        tagVMem_176 <= _GEN_690;
      end
    end else begin
      tagVMem_176 <= _GEN_690;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_177 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_177 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_177 <= _GEN_965;
      end else begin
        tagVMem_177 <= _GEN_691;
      end
    end else begin
      tagVMem_177 <= _GEN_691;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_178 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_178 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_178 <= _GEN_966;
      end else begin
        tagVMem_178 <= _GEN_692;
      end
    end else begin
      tagVMem_178 <= _GEN_692;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_179 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_179 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_179 <= _GEN_967;
      end else begin
        tagVMem_179 <= _GEN_693;
      end
    end else begin
      tagVMem_179 <= _GEN_693;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_180 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_180 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_180 <= _GEN_968;
      end else begin
        tagVMem_180 <= _GEN_694;
      end
    end else begin
      tagVMem_180 <= _GEN_694;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_181 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_181 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_181 <= _GEN_969;
      end else begin
        tagVMem_181 <= _GEN_695;
      end
    end else begin
      tagVMem_181 <= _GEN_695;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_182 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_182 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_182 <= _GEN_970;
      end else begin
        tagVMem_182 <= _GEN_696;
      end
    end else begin
      tagVMem_182 <= _GEN_696;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_183 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_183 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_183 <= _GEN_971;
      end else begin
        tagVMem_183 <= _GEN_697;
      end
    end else begin
      tagVMem_183 <= _GEN_697;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_184 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_184 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_184 <= _GEN_972;
      end else begin
        tagVMem_184 <= _GEN_698;
      end
    end else begin
      tagVMem_184 <= _GEN_698;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_185 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_185 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_185 <= _GEN_973;
      end else begin
        tagVMem_185 <= _GEN_699;
      end
    end else begin
      tagVMem_185 <= _GEN_699;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_186 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_186 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_186 <= _GEN_974;
      end else begin
        tagVMem_186 <= _GEN_700;
      end
    end else begin
      tagVMem_186 <= _GEN_700;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_187 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_187 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_187 <= _GEN_975;
      end else begin
        tagVMem_187 <= _GEN_701;
      end
    end else begin
      tagVMem_187 <= _GEN_701;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_188 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_188 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_188 <= _GEN_976;
      end else begin
        tagVMem_188 <= _GEN_702;
      end
    end else begin
      tagVMem_188 <= _GEN_702;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_189 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_189 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_189 <= _GEN_977;
      end else begin
        tagVMem_189 <= _GEN_703;
      end
    end else begin
      tagVMem_189 <= _GEN_703;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_190 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_190 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_190 <= _GEN_978;
      end else begin
        tagVMem_190 <= _GEN_704;
      end
    end else begin
      tagVMem_190 <= _GEN_704;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_191 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_191 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_191 <= _GEN_979;
      end else begin
        tagVMem_191 <= _GEN_705;
      end
    end else begin
      tagVMem_191 <= _GEN_705;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_192 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_192 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_192 <= _GEN_980;
      end else begin
        tagVMem_192 <= _GEN_706;
      end
    end else begin
      tagVMem_192 <= _GEN_706;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_193 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_193 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_193 <= _GEN_981;
      end else begin
        tagVMem_193 <= _GEN_707;
      end
    end else begin
      tagVMem_193 <= _GEN_707;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_194 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_194 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_194 <= _GEN_982;
      end else begin
        tagVMem_194 <= _GEN_708;
      end
    end else begin
      tagVMem_194 <= _GEN_708;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_195 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_195 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_195 <= _GEN_983;
      end else begin
        tagVMem_195 <= _GEN_709;
      end
    end else begin
      tagVMem_195 <= _GEN_709;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_196 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_196 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_196 <= _GEN_984;
      end else begin
        tagVMem_196 <= _GEN_710;
      end
    end else begin
      tagVMem_196 <= _GEN_710;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_197 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_197 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_197 <= _GEN_985;
      end else begin
        tagVMem_197 <= _GEN_711;
      end
    end else begin
      tagVMem_197 <= _GEN_711;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_198 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_198 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_198 <= _GEN_986;
      end else begin
        tagVMem_198 <= _GEN_712;
      end
    end else begin
      tagVMem_198 <= _GEN_712;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_199 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_199 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_199 <= _GEN_987;
      end else begin
        tagVMem_199 <= _GEN_713;
      end
    end else begin
      tagVMem_199 <= _GEN_713;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_200 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_200 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_200 <= _GEN_988;
      end else begin
        tagVMem_200 <= _GEN_714;
      end
    end else begin
      tagVMem_200 <= _GEN_714;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_201 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_201 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_201 <= _GEN_989;
      end else begin
        tagVMem_201 <= _GEN_715;
      end
    end else begin
      tagVMem_201 <= _GEN_715;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_202 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_202 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_202 <= _GEN_990;
      end else begin
        tagVMem_202 <= _GEN_716;
      end
    end else begin
      tagVMem_202 <= _GEN_716;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_203 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_203 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_203 <= _GEN_991;
      end else begin
        tagVMem_203 <= _GEN_717;
      end
    end else begin
      tagVMem_203 <= _GEN_717;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_204 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_204 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_204 <= _GEN_992;
      end else begin
        tagVMem_204 <= _GEN_718;
      end
    end else begin
      tagVMem_204 <= _GEN_718;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_205 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_205 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_205 <= _GEN_993;
      end else begin
        tagVMem_205 <= _GEN_719;
      end
    end else begin
      tagVMem_205 <= _GEN_719;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_206 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_206 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_206 <= _GEN_994;
      end else begin
        tagVMem_206 <= _GEN_720;
      end
    end else begin
      tagVMem_206 <= _GEN_720;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_207 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_207 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_207 <= _GEN_995;
      end else begin
        tagVMem_207 <= _GEN_721;
      end
    end else begin
      tagVMem_207 <= _GEN_721;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_208 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_208 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_208 <= _GEN_996;
      end else begin
        tagVMem_208 <= _GEN_722;
      end
    end else begin
      tagVMem_208 <= _GEN_722;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_209 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_209 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_209 <= _GEN_997;
      end else begin
        tagVMem_209 <= _GEN_723;
      end
    end else begin
      tagVMem_209 <= _GEN_723;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_210 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_210 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_210 <= _GEN_998;
      end else begin
        tagVMem_210 <= _GEN_724;
      end
    end else begin
      tagVMem_210 <= _GEN_724;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_211 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_211 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_211 <= _GEN_999;
      end else begin
        tagVMem_211 <= _GEN_725;
      end
    end else begin
      tagVMem_211 <= _GEN_725;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_212 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_212 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_212 <= _GEN_1000;
      end else begin
        tagVMem_212 <= _GEN_726;
      end
    end else begin
      tagVMem_212 <= _GEN_726;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_213 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_213 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_213 <= _GEN_1001;
      end else begin
        tagVMem_213 <= _GEN_727;
      end
    end else begin
      tagVMem_213 <= _GEN_727;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_214 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_214 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_214 <= _GEN_1002;
      end else begin
        tagVMem_214 <= _GEN_728;
      end
    end else begin
      tagVMem_214 <= _GEN_728;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_215 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_215 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_215 <= _GEN_1003;
      end else begin
        tagVMem_215 <= _GEN_729;
      end
    end else begin
      tagVMem_215 <= _GEN_729;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_216 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_216 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_216 <= _GEN_1004;
      end else begin
        tagVMem_216 <= _GEN_730;
      end
    end else begin
      tagVMem_216 <= _GEN_730;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_217 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_217 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_217 <= _GEN_1005;
      end else begin
        tagVMem_217 <= _GEN_731;
      end
    end else begin
      tagVMem_217 <= _GEN_731;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_218 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_218 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_218 <= _GEN_1006;
      end else begin
        tagVMem_218 <= _GEN_732;
      end
    end else begin
      tagVMem_218 <= _GEN_732;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_219 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_219 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_219 <= _GEN_1007;
      end else begin
        tagVMem_219 <= _GEN_733;
      end
    end else begin
      tagVMem_219 <= _GEN_733;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_220 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_220 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_220 <= _GEN_1008;
      end else begin
        tagVMem_220 <= _GEN_734;
      end
    end else begin
      tagVMem_220 <= _GEN_734;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_221 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_221 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_221 <= _GEN_1009;
      end else begin
        tagVMem_221 <= _GEN_735;
      end
    end else begin
      tagVMem_221 <= _GEN_735;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_222 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_222 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_222 <= _GEN_1010;
      end else begin
        tagVMem_222 <= _GEN_736;
      end
    end else begin
      tagVMem_222 <= _GEN_736;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_223 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_223 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_223 <= _GEN_1011;
      end else begin
        tagVMem_223 <= _GEN_737;
      end
    end else begin
      tagVMem_223 <= _GEN_737;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_224 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_224 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_224 <= _GEN_1012;
      end else begin
        tagVMem_224 <= _GEN_738;
      end
    end else begin
      tagVMem_224 <= _GEN_738;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_225 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_225 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_225 <= _GEN_1013;
      end else begin
        tagVMem_225 <= _GEN_739;
      end
    end else begin
      tagVMem_225 <= _GEN_739;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_226 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_226 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_226 <= _GEN_1014;
      end else begin
        tagVMem_226 <= _GEN_740;
      end
    end else begin
      tagVMem_226 <= _GEN_740;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_227 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_227 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_227 <= _GEN_1015;
      end else begin
        tagVMem_227 <= _GEN_741;
      end
    end else begin
      tagVMem_227 <= _GEN_741;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_228 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_228 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_228 <= _GEN_1016;
      end else begin
        tagVMem_228 <= _GEN_742;
      end
    end else begin
      tagVMem_228 <= _GEN_742;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_229 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_229 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_229 <= _GEN_1017;
      end else begin
        tagVMem_229 <= _GEN_743;
      end
    end else begin
      tagVMem_229 <= _GEN_743;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_230 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_230 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_230 <= _GEN_1018;
      end else begin
        tagVMem_230 <= _GEN_744;
      end
    end else begin
      tagVMem_230 <= _GEN_744;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_231 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_231 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_231 <= _GEN_1019;
      end else begin
        tagVMem_231 <= _GEN_745;
      end
    end else begin
      tagVMem_231 <= _GEN_745;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_232 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_232 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_232 <= _GEN_1020;
      end else begin
        tagVMem_232 <= _GEN_746;
      end
    end else begin
      tagVMem_232 <= _GEN_746;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_233 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_233 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_233 <= _GEN_1021;
      end else begin
        tagVMem_233 <= _GEN_747;
      end
    end else begin
      tagVMem_233 <= _GEN_747;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_234 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_234 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_234 <= _GEN_1022;
      end else begin
        tagVMem_234 <= _GEN_748;
      end
    end else begin
      tagVMem_234 <= _GEN_748;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_235 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_235 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_235 <= _GEN_1023;
      end else begin
        tagVMem_235 <= _GEN_749;
      end
    end else begin
      tagVMem_235 <= _GEN_749;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_236 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_236 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_236 <= _GEN_1024;
      end else begin
        tagVMem_236 <= _GEN_750;
      end
    end else begin
      tagVMem_236 <= _GEN_750;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_237 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_237 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_237 <= _GEN_1025;
      end else begin
        tagVMem_237 <= _GEN_751;
      end
    end else begin
      tagVMem_237 <= _GEN_751;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_238 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_238 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_238 <= _GEN_1026;
      end else begin
        tagVMem_238 <= _GEN_752;
      end
    end else begin
      tagVMem_238 <= _GEN_752;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_239 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_239 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_239 <= _GEN_1027;
      end else begin
        tagVMem_239 <= _GEN_753;
      end
    end else begin
      tagVMem_239 <= _GEN_753;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_240 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_240 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_240 <= _GEN_1028;
      end else begin
        tagVMem_240 <= _GEN_754;
      end
    end else begin
      tagVMem_240 <= _GEN_754;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_241 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_241 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_241 <= _GEN_1029;
      end else begin
        tagVMem_241 <= _GEN_755;
      end
    end else begin
      tagVMem_241 <= _GEN_755;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_242 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_242 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_242 <= _GEN_1030;
      end else begin
        tagVMem_242 <= _GEN_756;
      end
    end else begin
      tagVMem_242 <= _GEN_756;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_243 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_243 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_243 <= _GEN_1031;
      end else begin
        tagVMem_243 <= _GEN_757;
      end
    end else begin
      tagVMem_243 <= _GEN_757;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_244 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_244 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_244 <= _GEN_1032;
      end else begin
        tagVMem_244 <= _GEN_758;
      end
    end else begin
      tagVMem_244 <= _GEN_758;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_245 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_245 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_245 <= _GEN_1033;
      end else begin
        tagVMem_245 <= _GEN_759;
      end
    end else begin
      tagVMem_245 <= _GEN_759;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_246 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_246 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_246 <= _GEN_1034;
      end else begin
        tagVMem_246 <= _GEN_760;
      end
    end else begin
      tagVMem_246 <= _GEN_760;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_247 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_247 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_247 <= _GEN_1035;
      end else begin
        tagVMem_247 <= _GEN_761;
      end
    end else begin
      tagVMem_247 <= _GEN_761;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_248 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_248 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_248 <= _GEN_1036;
      end else begin
        tagVMem_248 <= _GEN_762;
      end
    end else begin
      tagVMem_248 <= _GEN_762;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_249 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_249 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_249 <= _GEN_1037;
      end else begin
        tagVMem_249 <= _GEN_763;
      end
    end else begin
      tagVMem_249 <= _GEN_763;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_250 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_250 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_250 <= _GEN_1038;
      end else begin
        tagVMem_250 <= _GEN_764;
      end
    end else begin
      tagVMem_250 <= _GEN_764;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_251 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_251 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_251 <= _GEN_1039;
      end else begin
        tagVMem_251 <= _GEN_765;
      end
    end else begin
      tagVMem_251 <= _GEN_765;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_252 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_252 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_252 <= _GEN_1040;
      end else begin
        tagVMem_252 <= _GEN_766;
      end
    end else begin
      tagVMem_252 <= _GEN_766;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_253 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_253 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_253 <= _GEN_1041;
      end else begin
        tagVMem_253 <= _GEN_767;
      end
    end else begin
      tagVMem_253 <= _GEN_767;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_254 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_254 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_254 <= _GEN_1042;
      end else begin
        tagVMem_254 <= _GEN_768;
      end
    end else begin
      tagVMem_254 <= _GEN_768;
    end
    if (reset) begin // @[DirectMappedCache.scala 42:24]
      tagVMem_255 <= 1'h0; // @[DirectMappedCache.scala 42:24]
    end else if (io_invalidate) begin // @[DirectMappedCache.scala 156:24]
      tagVMem_255 <= 1'h0; // @[DirectMappedCache.scala 157:19]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp == 2'h3) begin // @[DirectMappedCache.scala 144:43]
        tagVMem_255 <= _GEN_1043;
      end else begin
        tagVMem_255 <= _GEN_769;
      end
    end else begin
      tagVMem_255 <= _GEN_769;
    end
    if (8'hff == io_master_M_Addr[11:4]) begin // @[DirectMappedCache.scala 49:17]
      tagV <= tagVMem_255; // @[DirectMappedCache.scala 49:17]
    end else if (8'hfe == io_master_M_Addr[11:4]) begin // @[DirectMappedCache.scala 49:17]
      tagV <= tagVMem_254; // @[DirectMappedCache.scala 49:17]
    end else if (8'hfd == io_master_M_Addr[11:4]) begin // @[DirectMappedCache.scala 49:17]
      tagV <= tagVMem_253; // @[DirectMappedCache.scala 49:17]
    end else if (8'hfc == io_master_M_Addr[11:4]) begin // @[DirectMappedCache.scala 49:17]
      tagV <= tagVMem_252; // @[DirectMappedCache.scala 49:17]
    end else begin
      tagV <= _GEN_251;
    end
    fillReg <= stateReg == 2'h2 & _T_49; // @[DirectMappedCache.scala 130:27 DirectMappedCache.scala 93:11]
    if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      wrAddrReg <= _T_48; // @[DirectMappedCache.scala 131:15]
    end else begin
      wrAddrReg <= io_master_M_Addr[11:2]; // @[DirectMappedCache.scala 57:13]
    end
    if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp != 2'h0) begin // @[DirectMappedCache.scala 133:44]
        wrDataReg <= io_slave_S_Data; // @[DirectMappedCache.scala 135:17]
      end else begin
        wrDataReg <= io_master_M_Data; // @[DirectMappedCache.scala 58:13]
      end
    end else begin
      wrDataReg <= io_master_M_Data; // @[DirectMappedCache.scala 58:13]
    end
    if (reset) begin // @[DirectMappedCache.scala 77:21]
      stateReg <= 2'h0; // @[DirectMappedCache.scala 77:21]
    end else if (stateReg == 2'h3) begin // @[DirectMappedCache.scala 150:30]
      stateReg <= 2'h0; // @[DirectMappedCache.scala 152:14]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp != 2'h0) begin // @[DirectMappedCache.scala 133:44]
        stateReg <= _GEN_781;
      end else begin
        stateReg <= _GEN_777;
      end
    end else begin
      stateReg <= _GEN_777;
    end
    if (reset) begin // @[DirectMappedCache.scala 79:24]
      burstCntReg <= 2'h0; // @[DirectMappedCache.scala 79:24]
    end else if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp != 2'h0) begin // @[DirectMappedCache.scala 133:44]
        burstCntReg <= _lo_T_1; // @[DirectMappedCache.scala 142:19]
      end
    end
    if (~tagValid & _T_28) begin // @[DirectMappedCache.scala 101:50]
      missIndexReg <= masterReg_Addr[3:2]; // @[DirectMappedCache.scala 103:18]
    end
    if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp != 2'h0) begin // @[DirectMappedCache.scala 133:44]
        if (burstCntReg == missIndexReg) begin // @[DirectMappedCache.scala 136:42]
          slaveReg_Resp <= io_slave_S_Resp; // @[DirectMappedCache.scala 137:18]
        end
      end
    end
    if (stateReg == 2'h2) begin // @[DirectMappedCache.scala 130:27]
      if (io_slave_S_Resp != 2'h0) begin // @[DirectMappedCache.scala 133:44]
        if (burstCntReg == missIndexReg) begin // @[DirectMappedCache.scala 136:42]
          slaveReg_Data <= io_slave_S_Data; // @[DirectMappedCache.scala 137:18]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  masterReg_Cmd = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  masterReg_Addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  masterReg_ByteEn = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  tagVMem_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  tagVMem_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  tagVMem_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  tagVMem_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  tagVMem_4 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  tagVMem_5 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  tagVMem_6 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  tagVMem_7 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  tagVMem_8 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  tagVMem_9 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  tagVMem_10 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  tagVMem_11 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  tagVMem_12 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  tagVMem_13 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  tagVMem_14 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  tagVMem_15 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  tagVMem_16 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  tagVMem_17 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  tagVMem_18 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  tagVMem_19 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  tagVMem_20 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  tagVMem_21 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  tagVMem_22 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  tagVMem_23 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  tagVMem_24 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  tagVMem_25 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  tagVMem_26 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  tagVMem_27 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  tagVMem_28 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  tagVMem_29 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  tagVMem_30 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  tagVMem_31 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  tagVMem_32 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  tagVMem_33 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  tagVMem_34 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  tagVMem_35 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  tagVMem_36 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  tagVMem_37 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  tagVMem_38 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  tagVMem_39 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  tagVMem_40 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  tagVMem_41 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  tagVMem_42 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  tagVMem_43 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  tagVMem_44 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  tagVMem_45 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  tagVMem_46 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  tagVMem_47 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  tagVMem_48 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  tagVMem_49 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  tagVMem_50 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  tagVMem_51 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  tagVMem_52 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  tagVMem_53 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  tagVMem_54 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  tagVMem_55 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  tagVMem_56 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  tagVMem_57 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  tagVMem_58 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  tagVMem_59 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  tagVMem_60 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  tagVMem_61 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tagVMem_62 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  tagVMem_63 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  tagVMem_64 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  tagVMem_65 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  tagVMem_66 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  tagVMem_67 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  tagVMem_68 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  tagVMem_69 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  tagVMem_70 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  tagVMem_71 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  tagVMem_72 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  tagVMem_73 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  tagVMem_74 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  tagVMem_75 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  tagVMem_76 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  tagVMem_77 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  tagVMem_78 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  tagVMem_79 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  tagVMem_80 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  tagVMem_81 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  tagVMem_82 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  tagVMem_83 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  tagVMem_84 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  tagVMem_85 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  tagVMem_86 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  tagVMem_87 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  tagVMem_88 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  tagVMem_89 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  tagVMem_90 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  tagVMem_91 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  tagVMem_92 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  tagVMem_93 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  tagVMem_94 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  tagVMem_95 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  tagVMem_96 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  tagVMem_97 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  tagVMem_98 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  tagVMem_99 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  tagVMem_100 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  tagVMem_101 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  tagVMem_102 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  tagVMem_103 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  tagVMem_104 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  tagVMem_105 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  tagVMem_106 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  tagVMem_107 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  tagVMem_108 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  tagVMem_109 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  tagVMem_110 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  tagVMem_111 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  tagVMem_112 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  tagVMem_113 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  tagVMem_114 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  tagVMem_115 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  tagVMem_116 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  tagVMem_117 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  tagVMem_118 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  tagVMem_119 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  tagVMem_120 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  tagVMem_121 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  tagVMem_122 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  tagVMem_123 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  tagVMem_124 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  tagVMem_125 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  tagVMem_126 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  tagVMem_127 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  tagVMem_128 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  tagVMem_129 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  tagVMem_130 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  tagVMem_131 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  tagVMem_132 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  tagVMem_133 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  tagVMem_134 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  tagVMem_135 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  tagVMem_136 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  tagVMem_137 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  tagVMem_138 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  tagVMem_139 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  tagVMem_140 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  tagVMem_141 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  tagVMem_142 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  tagVMem_143 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  tagVMem_144 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  tagVMem_145 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  tagVMem_146 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  tagVMem_147 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  tagVMem_148 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  tagVMem_149 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  tagVMem_150 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  tagVMem_151 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  tagVMem_152 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  tagVMem_153 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tagVMem_154 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  tagVMem_155 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  tagVMem_156 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  tagVMem_157 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  tagVMem_158 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  tagVMem_159 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  tagVMem_160 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  tagVMem_161 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  tagVMem_162 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  tagVMem_163 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  tagVMem_164 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  tagVMem_165 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  tagVMem_166 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  tagVMem_167 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  tagVMem_168 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  tagVMem_169 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  tagVMem_170 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  tagVMem_171 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  tagVMem_172 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  tagVMem_173 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  tagVMem_174 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  tagVMem_175 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  tagVMem_176 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  tagVMem_177 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  tagVMem_178 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  tagVMem_179 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  tagVMem_180 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  tagVMem_181 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  tagVMem_182 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  tagVMem_183 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  tagVMem_184 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  tagVMem_185 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  tagVMem_186 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  tagVMem_187 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  tagVMem_188 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  tagVMem_189 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  tagVMem_190 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  tagVMem_191 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  tagVMem_192 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  tagVMem_193 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  tagVMem_194 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  tagVMem_195 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  tagVMem_196 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  tagVMem_197 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  tagVMem_198 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  tagVMem_199 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  tagVMem_200 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  tagVMem_201 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  tagVMem_202 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  tagVMem_203 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  tagVMem_204 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  tagVMem_205 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  tagVMem_206 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  tagVMem_207 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  tagVMem_208 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  tagVMem_209 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  tagVMem_210 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  tagVMem_211 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  tagVMem_212 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  tagVMem_213 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  tagVMem_214 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  tagVMem_215 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  tagVMem_216 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  tagVMem_217 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  tagVMem_218 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  tagVMem_219 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  tagVMem_220 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  tagVMem_221 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  tagVMem_222 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  tagVMem_223 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  tagVMem_224 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  tagVMem_225 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  tagVMem_226 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  tagVMem_227 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  tagVMem_228 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  tagVMem_229 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  tagVMem_230 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  tagVMem_231 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  tagVMem_232 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  tagVMem_233 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  tagVMem_234 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  tagVMem_235 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  tagVMem_236 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  tagVMem_237 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  tagVMem_238 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  tagVMem_239 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  tagVMem_240 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  tagVMem_241 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  tagVMem_242 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  tagVMem_243 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  tagVMem_244 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  tagVMem_245 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  tagVMem_246 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  tagVMem_247 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  tagVMem_248 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  tagVMem_249 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  tagVMem_250 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  tagVMem_251 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  tagVMem_252 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  tagVMem_253 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  tagVMem_254 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  tagVMem_255 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  tagV = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  fillReg = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  wrAddrReg = _RAND_261[9:0];
  _RAND_262 = {1{`RANDOM}};
  wrDataReg = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  stateReg = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  burstCntReg = _RAND_264[1:0];
  _RAND_265 = {1{`RANDOM}};
  missIndexReg = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  slaveReg_Resp = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  slaveReg_Data = _RAND_267[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemBlock_9(
  input        clock,
  input  [8:0] io_rdAddr,
  output [7:0] io_rdData,
  input  [8:0] io_wrAddr,
  input        io_wrEna,
  input  [7:0] io_wrData
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] mem [0:511];
  wire [7:0] mem_MPORT_1_data;
  wire [8:0] mem_MPORT_1_addr;
  wire [7:0] mem_MPORT_data;
  wire [8:0] mem_MPORT_addr;
  wire  mem_MPORT_mask;
  wire  mem_MPORT_en;
  reg [8:0] rdAddrReg; // @[MemBlock.scala 59:22]
  assign mem_MPORT_1_addr = rdAddrReg;
  assign mem_MPORT_1_data = mem[mem_MPORT_1_addr];
  assign mem_MPORT_data = io_wrData;
  assign mem_MPORT_addr = io_wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wrEna;
  assign io_rdData = mem_MPORT_1_data; // @[MemBlock.scala 60:13]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data;
    end
    rdAddrReg <= io_rdAddr; // @[MemBlock.scala 59:22]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rdAddrReg = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StackCache(
  input         clock,
  input         reset,
  input         io_ena_in,
  input  [2:0]  io_exsc_op,
  input  [31:0] io_exsc_opData,
  input  [31:0] io_exsc_opOff,
  output [31:0] io_scex_stackTop,
  output [31:0] io_scex_memTop,
  output        io_illMem,
  output        io_stall,
  input  [2:0]  io_fromCPU_M_Cmd,
  input  [31:0] io_fromCPU_M_Addr,
  input  [31:0] io_fromCPU_M_Data,
  input  [3:0]  io_fromCPU_M_ByteEn,
  output [1:0]  io_fromCPU_S_Resp,
  output [31:0] io_fromCPU_S_Data,
  output [2:0]  io_toMemory_M_Cmd,
  output [31:0] io_toMemory_M_Addr,
  output [31:0] io_toMemory_M_Data,
  output        io_toMemory_M_DataValid,
  output [3:0]  io_toMemory_M_DataByteEn,
  input  [1:0]  io_toMemory_S_Resp,
  input  [31:0] io_toMemory_S_Data,
  input         io_toMemory_S_CmdAccept
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  MemBlock_clock; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_io_rdData; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_io_wrData; // @[MemBlock.scala 15:11]
  wire  MemBlock_1_clock; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_1_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_1_io_rdData; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_1_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_1_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_1_io_wrData; // @[MemBlock.scala 15:11]
  wire  MemBlock_2_clock; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_2_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_2_io_rdData; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_2_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_2_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_2_io_wrData; // @[MemBlock.scala 15:11]
  wire  MemBlock_3_clock; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_3_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_3_io_rdData; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_3_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_3_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_3_io_wrData; // @[MemBlock.scala 15:11]
  reg [2:0] stateReg; // @[StackCache.scala 74:21]
  reg  isReserveReg; // @[StackCache.scala 77:25]
  reg [31:0] stackTopReg; // @[StackCache.scala 80:24]
  reg [31:0] memTopReg; // @[StackCache.scala 83:22]
  reg [32:0] transferAddrReg; // @[StackCache.scala 86:28]
  reg [31:0] newMemTopReg; // @[StackCache.scala 89:25]
  wire [23:0] _T_1 = {MemBlock_2_io_rdData,MemBlock_1_io_rdData,MemBlock_io_rdData}; // @[StackCache.scala 98:67]
  reg [8:0] rdAddrReg; // @[StackCache.scala 104:22]
  reg [1:0] responseToCPUReg; // @[StackCache.scala 107:29]
  wire [31:0] _T_3 = stackTopReg + 32'h800; // @[StackCache.scala 111:39]
  wire [32:0] _GEN_135 = {{1'd0}, _T_3}; // @[StackCache.scala 111:60]
  wire [32:0] _GEN_136 = {{1'd0}, memTopReg}; // @[StackCache.scala 111:100]
  wire  _T_5 = transferAddrReg < _GEN_136; // @[StackCache.scala 111:100]
  wire  _T_6 = _GEN_135 <= transferAddrReg & transferAddrReg < _GEN_136; // @[StackCache.scala 111:80]
  wire [32:0] _GEN_137 = {{1'd0}, newMemTopReg}; // @[StackCache.scala 112:39]
  wire  _T_7 = _GEN_137 <= transferAddrReg; // @[StackCache.scala 112:39]
  wire  _T_9 = _GEN_137 <= transferAddrReg & _T_5; // @[StackCache.scala 112:59]
  wire  writeEnable = isReserveReg ? _T_6 : _T_9; // @[StackCache.scala 110:24]
  wire [31:0] _T_14 = io_fromCPU_M_Addr + stackTopReg; // @[StackCache.scala 125:36]
  wire [8:0] relAddr = _T_14[10:2]; // @[StackCache.scala 125:50]
  wire [1:0] burstCounter = transferAddrReg[3:2]; // @[StackCache.scala 136:37]
  wire [31:0] stackTopInc = stackTopReg + io_exsc_opOff; // @[StackCache.scala 141:33]
  wire [31:0] _T_17 = memTopReg - stackTopReg; // @[StackCache.scala 142:33]
  wire  stackAboveMem = _T_17 < io_exsc_opOff; // @[StackCache.scala 142:47]
  wire  _T_18 = 3'h0 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_19 = 3'h0 == io_exsc_op; // @[Conditional.scala 37:30]
  wire  _T_20 = 3'h1 == io_exsc_op; // @[Conditional.scala 37:30]
  wire  _T_21 = 3'h2 == io_exsc_op; // @[Conditional.scala 37:30]
  wire  _T_22 = 3'h4 == io_exsc_op; // @[Conditional.scala 37:30]
  wire [31:0] _T_25 = {memTopReg[31:4],4'h0}; // @[StackCache.scala 166:67]
  wire [2:0] _T_26 = stackAboveMem ? 3'h1 : 3'h0; // @[StackCache.scala 172:26]
  wire  _T_27 = 3'h5 == io_exsc_op; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_0 = stackAboveMem ? stackTopInc : memTopReg; // @[StackCache.scala 178:31 StackCache.scala 179:23 StackCache.scala 83:22]
  wire  _T_28 = 3'h3 == io_exsc_op; // @[Conditional.scala 37:30]
  wire [31:0] _T_30 = stackTopReg - io_exsc_opOff; // @[StackCache.scala 186:42]
  wire [31:0] _T_32 = _T_30 + 32'h800; // @[StackCache.scala 190:27]
  wire [31:0] _T_35 = {_T_32[31:4],4'h0}; // @[StackCache.scala 190:73]
  wire [31:0] _T_38 = memTopReg - _T_30; // @[StackCache.scala 196:39]
  wire  _T_39 = _T_38 > 32'h800; // @[StackCache.scala 196:55]
  wire [2:0] _T_40 = _T_39 ? 3'h4 : 3'h0; // @[StackCache.scala 197:26]
  wire  _T_41 = 3'h6 == io_exsc_op; // @[Conditional.scala 37:30]
  wire [31:0] _T_43 = memTopReg - io_exsc_opOff; // @[StackCache.scala 203:41]
  wire [31:0] _T_46 = {_T_43[31:4],4'h0}; // @[StackCache.scala 205:52]
  wire  _GEN_1 = _T_41 ? 1'h0 : isReserveReg; // @[Conditional.scala 39:67 StackCache.scala 201:24 StackCache.scala 77:25]
  wire [8:0] _GEN_2 = _T_41 ? _T_46[10:2] : relAddr; // @[Conditional.scala 39:67 StackCache.scala 207:21 StackCache.scala 126:13]
  wire [32:0] _GEN_3 = _T_41 ? {{1'd0}, _T_46} : transferAddrReg; // @[Conditional.scala 39:67 StackCache.scala 209:27 StackCache.scala 86:28]
  wire [31:0] _GEN_4 = _T_41 ? _T_43 : newMemTopReg; // @[Conditional.scala 39:67 StackCache.scala 211:24 StackCache.scala 89:25]
  wire [2:0] _GEN_5 = _T_41 ? 3'h4 : 3'h0; // @[Conditional.scala 39:67 StackCache.scala 213:20 StackCache.scala 150:16]
  wire  _GEN_6 = _T_28 | _GEN_1; // @[Conditional.scala 39:67 StackCache.scala 184:24]
  wire [31:0] _GEN_7 = _T_28 ? _T_30 : stackTopReg; // @[Conditional.scala 39:67 StackCache.scala 187:23 StackCache.scala 80:24]
  wire [8:0] _GEN_8 = _T_28 ? _T_35[10:2] : _GEN_2; // @[Conditional.scala 39:67 StackCache.scala 192:21]
  wire [32:0] _GEN_9 = _T_28 ? {{1'd0}, _T_35} : _GEN_3; // @[Conditional.scala 39:67 StackCache.scala 194:27]
  wire [2:0] _GEN_10 = _T_28 ? _T_40 : _GEN_5; // @[Conditional.scala 39:67 StackCache.scala 197:20]
  wire [31:0] _GEN_11 = _T_28 ? newMemTopReg : _GEN_4; // @[Conditional.scala 39:67 StackCache.scala 89:25]
  wire [31:0] _GEN_12 = _T_27 ? stackTopInc : _GEN_7; // @[Conditional.scala 39:67 StackCache.scala 176:23]
  wire [31:0] _GEN_13 = _T_27 ? _GEN_0 : memTopReg; // @[Conditional.scala 39:67 StackCache.scala 83:22]
  wire  _GEN_14 = _T_27 ? isReserveReg : _GEN_6; // @[Conditional.scala 39:67 StackCache.scala 77:25]
  wire [8:0] _GEN_15 = _T_27 ? relAddr : _GEN_8; // @[Conditional.scala 39:67 StackCache.scala 126:13]
  wire [32:0] _GEN_16 = _T_27 ? transferAddrReg : _GEN_9; // @[Conditional.scala 39:67 StackCache.scala 86:28]
  wire [2:0] _GEN_17 = _T_27 ? 3'h0 : _GEN_10; // @[Conditional.scala 39:67 StackCache.scala 150:16]
  wire [31:0] _GEN_18 = _T_27 ? newMemTopReg : _GEN_11; // @[Conditional.scala 39:67 StackCache.scala 89:25]
  wire [32:0] _GEN_19 = _T_22 ? {{1'd0}, _T_25} : _GEN_16; // @[Conditional.scala 39:67 StackCache.scala 166:27]
  wire [31:0] _GEN_20 = _T_22 ? stackTopInc : _GEN_18; // @[Conditional.scala 39:67 StackCache.scala 169:24]
  wire [2:0] _GEN_21 = _T_22 ? _T_26 : _GEN_17; // @[Conditional.scala 39:67 StackCache.scala 172:20]
  wire [31:0] _GEN_22 = _T_22 ? stackTopReg : _GEN_12; // @[Conditional.scala 39:67 StackCache.scala 80:24]
  wire [31:0] _GEN_23 = _T_22 ? memTopReg : _GEN_13; // @[Conditional.scala 39:67 StackCache.scala 83:22]
  wire  _GEN_24 = _T_22 ? isReserveReg : _GEN_14; // @[Conditional.scala 39:67 StackCache.scala 77:25]
  wire [8:0] _GEN_25 = _T_22 ? relAddr : _GEN_15; // @[Conditional.scala 39:67 StackCache.scala 126:13]
  wire [31:0] _GEN_26 = _T_21 ? io_exsc_opData : _GEN_23; // @[Conditional.scala 39:67 StackCache.scala 162:21]
  wire [32:0] _GEN_27 = _T_21 ? transferAddrReg : _GEN_19; // @[Conditional.scala 39:67 StackCache.scala 86:28]
  wire [2:0] _GEN_29 = _T_21 ? 3'h0 : _GEN_21; // @[Conditional.scala 39:67 StackCache.scala 150:16]
  wire [31:0] _GEN_30 = _T_21 ? stackTopReg : _GEN_22; // @[Conditional.scala 39:67 StackCache.scala 80:24]
  wire [8:0] _GEN_32 = _T_21 ? relAddr : _GEN_25; // @[Conditional.scala 39:67 StackCache.scala 126:13]
  wire [2:0] _GEN_37 = _T_20 ? 3'h0 : _GEN_29; // @[Conditional.scala 39:67 StackCache.scala 150:16]
  wire [8:0] _GEN_39 = _T_20 ? relAddr : _GEN_32; // @[Conditional.scala 39:67 StackCache.scala 126:13]
  wire [8:0] _GEN_46 = _T_19 ? relAddr : _GEN_39; // @[Conditional.scala 40:58 StackCache.scala 126:13]
  wire  _T_48 = 3'h4 == stateReg; // @[Conditional.scala 37:30]
  wire [32:0] _T_50 = transferAddrReg + 33'h4; // @[StackCache.scala 222:46]
  wire [8:0] _T_53 = io_toMemory_S_CmdAccept ? _T_50[10:2] : rdAddrReg; // @[StackCache.scala 232:23]
  wire [2:0] _T_55 = io_toMemory_S_CmdAccept ? 3'h3 : 3'h4; // @[StackCache.scala 238:22]
  wire  _T_56 = 3'h3 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_60 = burstCounter == 2'h3; // @[StackCache.scala 257:36]
  wire [2:0] _T_61 = burstCounter == 2'h3 ? 3'h5 : 3'h3; // @[StackCache.scala 257:22]
  wire  _T_62 = 3'h5 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_63 = _GEN_136 <= transferAddrReg; // @[StackCache.scala 263:36]
  wire  _T_64 = io_toMemory_S_Resp == 2'h1; // @[StackCache.scala 267:42]
  wire [2:0] _T_65 = _T_63 ? 3'h0 : 3'h4; // @[StackCache.scala 268:26]
  wire  _T_66 = io_toMemory_S_Resp == 2'h3; // @[StackCache.scala 269:46]
  wire [2:0] _T_67 = io_toMemory_S_Resp == 2'h3 ? 3'h0 : 3'h5; // @[StackCache.scala 269:26]
  wire [2:0] _T_68 = io_toMemory_S_Resp == 2'h1 ? _T_65 : _T_67; // @[StackCache.scala 267:22]
  wire [31:0] _T_72 = isReserveReg ? _T_3 : newMemTopReg; // @[StackCache.scala 275:27]
  wire [31:0] _T_73 = _T_63 ? _T_72 : memTopReg; // @[StackCache.scala 274:23]
  wire  _T_74 = 3'h1 == stateReg; // @[Conditional.scala 37:30]
  wire [2:0] _T_76 = io_toMemory_S_CmdAccept ? 3'h2 : 3'h1; // @[StackCache.scala 295:22]
  wire  _T_77 = 3'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _T_82 = ~_T_7 & _T_63; // @[StackCache.scala 309:40]
  wire [3:0] _T_84 = _T_82 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_89 = _T_7 ? 3'h0 : 3'h1; // @[StackCache.scala 321:14]
  wire [2:0] _T_90 = _T_60 ? _T_89 : 3'h2; // @[StackCache.scala 320:24]
  wire [31:0] _T_91 = _T_7 ? newMemTopReg : memTopReg; // @[StackCache.scala 325:25]
  wire [3:0] _GEN_49 = _T_64 ? _T_84 : 4'h0; // @[StackCache.scala 304:48 StackCache.scala 312:18 StackCache.scala 128:13]
  wire [31:0] _GEN_50 = _T_64 ? io_toMemory_S_Data : io_fromCPU_M_Data; // @[StackCache.scala 304:48 StackCache.scala 313:19 StackCache.scala 129:13]
  wire [8:0] _GEN_51 = _T_64 ? transferAddrReg[10:2] : relAddr; // @[StackCache.scala 304:48 StackCache.scala 314:19 StackCache.scala 127:13]
  wire [32:0] _GEN_52 = _T_64 ? _T_50 : transferAddrReg; // @[StackCache.scala 304:48 StackCache.scala 317:25 StackCache.scala 86:28]
  wire [2:0] _GEN_53 = _T_64 ? _T_90 : stateReg; // @[StackCache.scala 304:48 StackCache.scala 320:18 StackCache.scala 74:21]
  wire [31:0] _GEN_54 = _T_64 ? _T_91 : memTopReg; // @[StackCache.scala 304:48 StackCache.scala 325:19 StackCache.scala 83:22]
  wire [32:0] _GEN_55 = _T_66 ? _T_50 : _GEN_52; // @[StackCache.scala 329:49 StackCache.scala 330:25]
  wire [2:0] _GEN_56 = _T_66 ? 3'h6 : _GEN_53; // @[StackCache.scala 329:49 StackCache.scala 331:18]
  wire  _T_95 = 3'h6 == stateReg; // @[Conditional.scala 37:30]
  wire [32:0] _GEN_57 = io_toMemory_S_Resp != 2'h0 ? _T_50 : transferAddrReg; // @[StackCache.scala 337:50 StackCache.scala 338:25 StackCache.scala 86:28]
  wire [2:0] _GEN_59 = _T_60 ? 3'h0 : stateReg; // @[StackCache.scala 340:54 StackCache.scala 342:18 StackCache.scala 74:21]
  wire [32:0] _GEN_60 = _T_95 ? _GEN_57 : transferAddrReg; // @[Conditional.scala 39:67 StackCache.scala 86:28]
  wire [2:0] _GEN_62 = _T_95 ? _GEN_59 : stateReg; // @[Conditional.scala 39:67 StackCache.scala 74:21]
  wire [3:0] _GEN_63 = _T_77 ? _GEN_49 : 4'h0; // @[Conditional.scala 39:67 StackCache.scala 128:13]
  wire [31:0] _GEN_64 = _T_77 ? _GEN_50 : io_fromCPU_M_Data; // @[Conditional.scala 39:67 StackCache.scala 129:13]
  wire [8:0] _GEN_65 = _T_77 ? _GEN_51 : relAddr; // @[Conditional.scala 39:67 StackCache.scala 127:13]
  wire [32:0] _GEN_66 = _T_77 ? _GEN_55 : _GEN_60; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_67 = _T_77 ? _GEN_56 : _GEN_62; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_68 = _T_77 ? _GEN_54 : memTopReg; // @[Conditional.scala 39:67 StackCache.scala 83:22]
  wire  _GEN_69 = _T_77 ? 1'h0 : _T_95 & _T_60; // @[Conditional.scala 39:67 StackCache.scala 115:13]
  wire [2:0] _GEN_70 = _T_74 ? 3'h2 : 3'h0; // @[Conditional.scala 39:67 StackCache.scala 289:25 StackCache.scala 118:21]
  wire [2:0] _GEN_71 = _T_74 ? _T_76 : _GEN_67; // @[Conditional.scala 39:67 StackCache.scala 295:16]
  wire [3:0] _GEN_73 = _T_74 ? 4'h0 : _GEN_63; // @[Conditional.scala 39:67 StackCache.scala 128:13]
  wire [31:0] _GEN_74 = _T_74 ? io_fromCPU_M_Data : _GEN_64; // @[Conditional.scala 39:67 StackCache.scala 129:13]
  wire [8:0] _GEN_75 = _T_74 ? relAddr : _GEN_65; // @[Conditional.scala 39:67 StackCache.scala 127:13]
  wire [32:0] _GEN_76 = _T_74 ? transferAddrReg : _GEN_66; // @[Conditional.scala 39:67 StackCache.scala 86:28]
  wire [31:0] _GEN_77 = _T_74 ? memTopReg : _GEN_68; // @[Conditional.scala 39:67 StackCache.scala 83:22]
  wire  _GEN_78 = _T_74 ? 1'h0 : _GEN_69; // @[Conditional.scala 39:67 StackCache.scala 115:13]
  wire [2:0] _GEN_79 = _T_62 ? _T_68 : _GEN_71; // @[Conditional.scala 39:67 StackCache.scala 267:16]
  wire  _GEN_80 = _T_62 ? _T_66 : _GEN_78; // @[Conditional.scala 39:67 StackCache.scala 271:17]
  wire [31:0] _GEN_81 = _T_62 ? _T_73 : _GEN_77; // @[Conditional.scala 39:67 StackCache.scala 274:17]
  wire [8:0] _GEN_82 = _T_62 ? rdAddrReg : relAddr; // @[Conditional.scala 39:67 StackCache.scala 281:17 StackCache.scala 126:13]
  wire [2:0] _GEN_83 = _T_62 ? 3'h0 : _GEN_70; // @[Conditional.scala 39:67 StackCache.scala 118:21]
  wire [3:0] _GEN_85 = _T_62 ? 4'h0 : _GEN_73; // @[Conditional.scala 39:67 StackCache.scala 128:13]
  wire [31:0] _GEN_86 = _T_62 ? io_fromCPU_M_Data : _GEN_74; // @[Conditional.scala 39:67 StackCache.scala 129:13]
  wire [8:0] _GEN_87 = _T_62 ? relAddr : _GEN_75; // @[Conditional.scala 39:67 StackCache.scala 127:13]
  wire [32:0] _GEN_88 = _T_62 ? transferAddrReg : _GEN_76; // @[Conditional.scala 39:67 StackCache.scala 86:28]
  wire [8:0] _GEN_89 = _T_56 ? _T_50[10:2] : _GEN_82; // @[Conditional.scala 39:67 StackCache.scala 249:17]
  wire [2:0] _GEN_92 = _T_56 ? _T_61 : _GEN_79; // @[Conditional.scala 39:67 StackCache.scala 257:16]
  wire  _GEN_93 = _T_56 ? 1'h0 : _GEN_80; // @[Conditional.scala 39:67 StackCache.scala 115:13]
  wire [2:0] _GEN_95 = _T_56 ? 3'h0 : _GEN_83; // @[Conditional.scala 39:67 StackCache.scala 118:21]
  wire [3:0] _GEN_97 = _T_56 ? 4'h0 : _GEN_85; // @[Conditional.scala 39:67 StackCache.scala 128:13]
  wire [31:0] _GEN_98 = _T_56 ? io_fromCPU_M_Data : _GEN_86; // @[Conditional.scala 39:67 StackCache.scala 129:13]
  wire [8:0] _GEN_99 = _T_56 ? relAddr : _GEN_87; // @[Conditional.scala 39:67 StackCache.scala 127:13]
  wire [2:0] _GEN_100 = _T_48 ? 3'h1 : _GEN_95; // @[Conditional.scala 39:67 StackCache.scala 225:25]
  wire  _GEN_101 = _T_48 | _T_56; // @[Conditional.scala 39:67 StackCache.scala 226:31]
  wire [8:0] _GEN_102 = _T_48 ? _T_53 : _GEN_89; // @[Conditional.scala 39:67 StackCache.scala 232:17]
  wire  _GEN_106 = _T_48 ? 1'h0 : _GEN_93; // @[Conditional.scala 39:67 StackCache.scala 115:13]
  wire [3:0] _GEN_109 = _T_48 ? 4'h0 : _GEN_97; // @[Conditional.scala 39:67 StackCache.scala 128:13]
  wire [31:0] _GEN_110 = _T_48 ? io_fromCPU_M_Data : _GEN_98; // @[Conditional.scala 39:67 StackCache.scala 129:13]
  wire [8:0] _GEN_111 = _T_48 ? relAddr : _GEN_99; // @[Conditional.scala 39:67 StackCache.scala 127:13]
  wire [2:0] _GEN_119 = _T_18 ? 3'h0 : _GEN_100; // @[Conditional.scala 40:58 StackCache.scala 118:21]
  wire [3:0] _GEN_124 = _T_18 ? 4'h0 : _GEN_109; // @[Conditional.scala 40:58 StackCache.scala 128:13]
  wire [31:0] mb_wrData = _T_18 ? io_fromCPU_M_Data : _GEN_110; // @[Conditional.scala 40:58 StackCache.scala 129:13]
  wire [3:0] mb_wrEna = io_fromCPU_M_Cmd == 3'h1 ? io_fromCPU_M_ByteEn : _GEN_124; // @[StackCache.scala 356:40 StackCache.scala 358:14]
  MemBlock_9 MemBlock ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_clock),
    .io_rdAddr(MemBlock_io_rdAddr),
    .io_rdData(MemBlock_io_rdData),
    .io_wrAddr(MemBlock_io_wrAddr),
    .io_wrEna(MemBlock_io_wrEna),
    .io_wrData(MemBlock_io_wrData)
  );
  MemBlock_9 MemBlock_1 ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_1_clock),
    .io_rdAddr(MemBlock_1_io_rdAddr),
    .io_rdData(MemBlock_1_io_rdData),
    .io_wrAddr(MemBlock_1_io_wrAddr),
    .io_wrEna(MemBlock_1_io_wrEna),
    .io_wrData(MemBlock_1_io_wrData)
  );
  MemBlock_9 MemBlock_2 ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_2_clock),
    .io_rdAddr(MemBlock_2_io_rdAddr),
    .io_rdData(MemBlock_2_io_rdData),
    .io_wrAddr(MemBlock_2_io_wrAddr),
    .io_wrEna(MemBlock_2_io_wrEna),
    .io_wrData(MemBlock_2_io_wrData)
  );
  MemBlock_9 MemBlock_3 ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_3_clock),
    .io_rdAddr(MemBlock_3_io_rdAddr),
    .io_rdData(MemBlock_3_io_rdData),
    .io_wrAddr(MemBlock_3_io_wrAddr),
    .io_wrEna(MemBlock_3_io_wrEna),
    .io_wrData(MemBlock_3_io_wrData)
  );
  assign io_scex_stackTop = stackTopReg; // @[StackCache.scala 132:20]
  assign io_scex_memTop = memTopReg; // @[StackCache.scala 133:18]
  assign io_illMem = _T_18 ? 1'h0 : _GEN_106; // @[Conditional.scala 40:58 StackCache.scala 115:13]
  assign io_stall = stateReg != 3'h0; // @[StackCache.scala 114:24]
  assign io_fromCPU_S_Resp = responseToCPUReg; // @[StackCache.scala 352:21]
  assign io_fromCPU_S_Data = {MemBlock_3_io_rdData,_T_1}; // @[StackCache.scala 98:67]
  assign io_toMemory_M_Cmd = ~io_ena_in ? 3'h0 : _GEN_119; // @[StackCache.scala 382:21 StackCache.scala 387:23]
  assign io_toMemory_M_Addr = transferAddrReg[31:0]; // @[StackCache.scala 119:22]
  assign io_toMemory_M_Data = {MemBlock_3_io_rdData,_T_1}; // @[StackCache.scala 98:67]
  assign io_toMemory_M_DataValid = _T_18 ? 1'h0 : _GEN_101; // @[Conditional.scala 40:58 StackCache.scala 121:27]
  assign io_toMemory_M_DataByteEn = writeEnable ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  assign MemBlock_clock = clock;
  assign MemBlock_io_rdAddr = _T_18 ? _GEN_46 : _GEN_102; // @[Conditional.scala 40:58]
  assign MemBlock_io_wrAddr = _T_18 ? relAddr : _GEN_111; // @[Conditional.scala 40:58 StackCache.scala 127:13]
  assign MemBlock_io_wrEna = mb_wrEna[0]; // @[StackCache.scala 373:32]
  assign MemBlock_io_wrData = mb_wrData[7:0]; // @[StackCache.scala 374:16]
  assign MemBlock_1_clock = clock;
  assign MemBlock_1_io_rdAddr = _T_18 ? _GEN_46 : _GEN_102; // @[Conditional.scala 40:58]
  assign MemBlock_1_io_wrAddr = _T_18 ? relAddr : _GEN_111; // @[Conditional.scala 40:58 StackCache.scala 127:13]
  assign MemBlock_1_io_wrEna = mb_wrEna[1]; // @[StackCache.scala 373:32]
  assign MemBlock_1_io_wrData = mb_wrData[15:8]; // @[StackCache.scala 374:16]
  assign MemBlock_2_clock = clock;
  assign MemBlock_2_io_rdAddr = _T_18 ? _GEN_46 : _GEN_102; // @[Conditional.scala 40:58]
  assign MemBlock_2_io_wrAddr = _T_18 ? relAddr : _GEN_111; // @[Conditional.scala 40:58 StackCache.scala 127:13]
  assign MemBlock_2_io_wrEna = mb_wrEna[2]; // @[StackCache.scala 373:32]
  assign MemBlock_2_io_wrData = mb_wrData[23:16]; // @[StackCache.scala 374:16]
  assign MemBlock_3_clock = clock;
  assign MemBlock_3_io_rdAddr = _T_18 ? _GEN_46 : _GEN_102; // @[Conditional.scala 40:58]
  assign MemBlock_3_io_wrAddr = _T_18 ? relAddr : _GEN_111; // @[Conditional.scala 40:58 StackCache.scala 127:13]
  assign MemBlock_3_io_wrEna = mb_wrEna[3]; // @[StackCache.scala 373:32]
  assign MemBlock_3_io_wrData = mb_wrData[31:24]; // @[StackCache.scala 374:16]
  always @(posedge clock) begin
    if (reset) begin // @[StackCache.scala 74:21]
      stateReg <= 3'h0; // @[StackCache.scala 74:21]
    end else if (!(~io_ena_in)) begin // @[StackCache.scala 382:21]
      if (_T_18) begin // @[Conditional.scala 40:58]
        if (_T_19) begin // @[Conditional.scala 40:58]
          stateReg <= 3'h0; // @[StackCache.scala 150:16]
        end else begin
          stateReg <= _GEN_37;
        end
      end else if (_T_48) begin // @[Conditional.scala 39:67]
        stateReg <= _T_55; // @[StackCache.scala 238:16]
      end else begin
        stateReg <= _GEN_92;
      end
    end
    if (_T_18) begin // @[Conditional.scala 40:58]
      if (!(_T_19)) begin // @[Conditional.scala 40:58]
        if (!(_T_20)) begin // @[Conditional.scala 39:67]
          if (!(_T_21)) begin // @[Conditional.scala 39:67]
            isReserveReg <= _GEN_24;
          end
        end
      end
    end
    if (!(~io_ena_in)) begin // @[StackCache.scala 382:21]
      if (_T_18) begin // @[Conditional.scala 40:58]
        if (!(_T_19)) begin // @[Conditional.scala 40:58]
          if (_T_20) begin // @[Conditional.scala 39:67]
            stackTopReg <= io_exsc_opData; // @[StackCache.scala 158:23]
          end else begin
            stackTopReg <= _GEN_30;
          end
        end
      end
    end
    if (!(~io_ena_in)) begin // @[StackCache.scala 382:21]
      if (_T_18) begin // @[Conditional.scala 40:58]
        if (!(_T_19)) begin // @[Conditional.scala 40:58]
          if (!(_T_20)) begin // @[Conditional.scala 39:67]
            memTopReg <= _GEN_26;
          end
        end
      end else if (!(_T_48)) begin // @[Conditional.scala 39:67]
        if (!(_T_56)) begin // @[Conditional.scala 39:67]
          memTopReg <= _GEN_81;
        end
      end
    end
    if (!(~io_ena_in)) begin // @[StackCache.scala 382:21]
      if (_T_18) begin // @[Conditional.scala 40:58]
        if (!(_T_19)) begin // @[Conditional.scala 40:58]
          if (!(_T_20)) begin // @[Conditional.scala 39:67]
            transferAddrReg <= _GEN_27;
          end
        end
      end else if (_T_48) begin // @[Conditional.scala 39:67]
        if (io_toMemory_S_CmdAccept) begin // @[StackCache.scala 235:29]
          transferAddrReg <= _T_50;
        end
      end else if (_T_56) begin // @[Conditional.scala 39:67]
        transferAddrReg <= _T_50; // @[StackCache.scala 255:23]
      end else begin
        transferAddrReg <= _GEN_88;
      end
    end
    if (_T_18) begin // @[Conditional.scala 40:58]
      if (!(_T_19)) begin // @[Conditional.scala 40:58]
        if (!(_T_20)) begin // @[Conditional.scala 39:67]
          if (!(_T_21)) begin // @[Conditional.scala 39:67]
            newMemTopReg <= _GEN_20;
          end
        end
      end
    end
    rdAddrReg <= MemBlock_io_rdAddr; // @[StackCache.scala 104:22]
    if (reset) begin // @[StackCache.scala 107:29]
      responseToCPUReg <= 2'h0; // @[StackCache.scala 107:29]
    end else if (io_fromCPU_M_Cmd == 3'h1) begin // @[StackCache.scala 356:40]
      responseToCPUReg <= 2'h1; // @[StackCache.scala 361:22]
    end else if (io_fromCPU_M_Cmd == 3'h2) begin // @[StackCache.scala 363:45]
      responseToCPUReg <= 2'h1; // @[StackCache.scala 365:22]
    end else begin
      responseToCPUReg <= 2'h0; // @[StackCache.scala 139:20]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  isReserveReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  stackTopReg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  memTopReg = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  transferAddrReg = _RAND_4[32:0];
  _RAND_5 = {1{`RANDOM}};
  newMemTopReg = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  rdAddrReg = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  responseToCPUReg = _RAND_7[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NullCache(
  input         clock,
  input         reset,
  input  [2:0]  io_master_M_Cmd,
  input  [31:0] io_master_M_Addr,
  output [1:0]  io_master_S_Resp,
  output [31:0] io_master_S_Data,
  output [2:0]  io_slave_M_Cmd,
  output [31:0] io_slave_M_Addr,
  input  [1:0]  io_slave_S_Resp,
  input  [31:0] io_slave_S_Data,
  input         io_slave_S_CmdAccept
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] stateReg; // @[NullCache.scala 32:21]
  reg [1:0] burstCntReg; // @[NullCache.scala 33:24]
  reg [1:0] posReg; // @[NullCache.scala 34:19]
  reg [2:0] masterReg_Cmd; // @[NullCache.scala 37:22]
  reg [31:0] masterReg_Addr; // @[NullCache.scala 37:22]
  reg [1:0] slaveReg_Resp; // @[NullCache.scala 40:21]
  reg [31:0] slaveReg_Data; // @[NullCache.scala 40:21]
  wire [27:0] hi = masterReg_Addr[31:4]; // @[NullCache.scala 51:40]
  wire [1:0] _GEN_7 = burstCntReg == 2'h3 ? 2'h2 : stateReg; // @[NullCache.scala 66:50 NullCache.scala 67:18 NullCache.scala 32:21]
  wire [1:0] _T_10 = burstCntReg + 2'h1; // @[NullCache.scala 69:34]
  wire [1:0] _GEN_8 = io_slave_S_Resp != 2'h0 ? _GEN_7 : stateReg; // @[NullCache.scala 65:44 NullCache.scala 32:21]
  wire [1:0] _GEN_12 = stateReg == 2'h1 ? _GEN_8 : stateReg; // @[NullCache.scala 61:27 NullCache.scala 32:21]
  wire [1:0] _GEN_16 = stateReg == 2'h2 ? 2'h0 : _GEN_12; // @[NullCache.scala 73:31 NullCache.scala 75:14]
  assign io_master_S_Resp = stateReg == 2'h2 ? slaveReg_Resp : 2'h0; // @[NullCache.scala 73:31 NullCache.scala 74:17 NullCache.scala 57:20]
  assign io_master_S_Data = stateReg == 2'h2 ? slaveReg_Data : 32'h0; // @[NullCache.scala 73:31 NullCache.scala 74:17 NullCache.scala 58:20]
  assign io_slave_M_Cmd = masterReg_Cmd == 3'h2 ? 3'h2 : 3'h0; // @[NullCache.scala 79:37 NullCache.scala 80:20 NullCache.scala 50:18]
  assign io_slave_M_Addr = {hi,4'h0}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (reset) begin // @[NullCache.scala 32:21]
      stateReg <= 2'h0; // @[NullCache.scala 32:21]
    end else if (masterReg_Cmd == 3'h2) begin // @[NullCache.scala 79:37]
      if (io_slave_S_CmdAccept) begin // @[NullCache.scala 81:44]
        stateReg <= 2'h1; // @[NullCache.scala 82:16]
      end else begin
        stateReg <= _GEN_16;
      end
    end else begin
      stateReg <= _GEN_16;
    end
    if (reset) begin // @[NullCache.scala 33:24]
      burstCntReg <= 2'h0; // @[NullCache.scala 33:24]
    end else if (stateReg == 2'h1) begin // @[NullCache.scala 61:27]
      if (io_slave_S_Resp != 2'h0) begin // @[NullCache.scala 65:44]
        burstCntReg <= _T_10; // @[NullCache.scala 69:19]
      end
    end
    if (masterReg_Cmd == 3'h2) begin // @[NullCache.scala 79:37]
      if (io_slave_S_CmdAccept) begin // @[NullCache.scala 81:44]
        posReg <= masterReg_Addr[3:2]; // @[NullCache.scala 83:14]
      end
    end
    if (reset) begin // @[NullCache.scala 45:15]
      masterReg_Cmd <= 3'h0; // @[NullCache.scala 46:19]
    end else if (masterReg_Cmd != 3'h2 | io_slave_S_CmdAccept) begin // @[NullCache.scala 42:73]
      masterReg_Cmd <= io_master_M_Cmd; // @[NullCache.scala 43:15]
    end
    if (masterReg_Cmd != 3'h2 | io_slave_S_CmdAccept) begin // @[NullCache.scala 42:73]
      masterReg_Addr <= io_master_M_Addr; // @[NullCache.scala 43:15]
    end
    if (stateReg == 2'h1) begin // @[NullCache.scala 61:27]
      if (burstCntReg == posReg) begin // @[NullCache.scala 62:34]
        slaveReg_Resp <= io_slave_S_Resp; // @[NullCache.scala 63:16]
      end
    end
    if (stateReg == 2'h1) begin // @[NullCache.scala 61:27]
      if (burstCntReg == posReg) begin // @[NullCache.scala 62:34]
        slaveReg_Data <= io_slave_S_Data; // @[NullCache.scala 63:16]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  burstCntReg = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  posReg = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  masterReg_Cmd = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  masterReg_Addr = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  slaveReg_Resp = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  slaveReg_Data = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module OcpBurstBus(
  output [2:0]  io_master_M_Cmd,
  output [31:0] io_master_M_Addr,
  output [31:0] io_master_M_Data,
  output        io_master_M_DataValid,
  output [3:0]  io_master_M_DataByteEn,
  input  [1:0]  io_master_S_Resp,
  input  [31:0] io_master_S_Data,
  input         io_master_S_CmdAccept,
  input         io_master_S_DataAccept,
  input  [2:0]  io_slave_M_Cmd,
  input  [31:0] io_slave_M_Addr,
  input  [31:0] io_slave_M_Data,
  input         io_slave_M_DataValid,
  input  [3:0]  io_slave_M_DataByteEn,
  output [1:0]  io_slave_S_Resp,
  output [31:0] io_slave_S_Data,
  output        io_slave_S_CmdAccept,
  output        io_slave_S_DataAccept
);
  assign io_master_M_Cmd = io_slave_M_Cmd; // @[OcpBurst.scala 244:15]
  assign io_master_M_Addr = io_slave_M_Addr; // @[OcpBurst.scala 244:15]
  assign io_master_M_Data = io_slave_M_Data; // @[OcpBurst.scala 244:15]
  assign io_master_M_DataValid = io_slave_M_DataValid; // @[OcpBurst.scala 244:15]
  assign io_master_M_DataByteEn = io_slave_M_DataByteEn; // @[OcpBurst.scala 244:15]
  assign io_slave_S_Resp = io_master_S_Resp; // @[OcpBurst.scala 245:14]
  assign io_slave_S_Data = io_master_S_Data; // @[OcpBurst.scala 245:14]
  assign io_slave_S_CmdAccept = io_master_S_CmdAccept; // @[OcpBurst.scala 245:14]
  assign io_slave_S_DataAccept = io_master_S_DataAccept; // @[OcpBurst.scala 245:14]
endmodule
module WriteNoBuffer(
  input         clock,
  input         reset,
  input  [2:0]  io_readMaster_M_Cmd,
  input  [31:0] io_readMaster_M_Addr,
  input  [31:0] io_readMaster_M_Data,
  input         io_readMaster_M_DataValid,
  input  [3:0]  io_readMaster_M_DataByteEn,
  output [1:0]  io_readMaster_S_Resp,
  output [31:0] io_readMaster_S_Data,
  output        io_readMaster_S_CmdAccept,
  output        io_readMaster_S_DataAccept,
  input  [2:0]  io_writeMaster_M_Cmd,
  input  [31:0] io_writeMaster_M_Addr,
  input  [31:0] io_writeMaster_M_Data,
  input  [3:0]  io_writeMaster_M_ByteEn,
  output [1:0]  io_writeMaster_S_Resp,
  output [2:0]  io_slave_M_Cmd,
  output [31:0] io_slave_M_Addr,
  output [31:0] io_slave_M_Data,
  output        io_slave_M_DataValid,
  output [3:0]  io_slave_M_DataByteEn,
  input  [1:0]  io_slave_S_Resp,
  input  [31:0] io_slave_S_Data,
  input         io_slave_S_CmdAccept,
  input         io_slave_S_DataAccept
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[WriteNoBuffer.scala 68:18]
  reg [1:0] cntReg; // @[WriteNoBuffer.scala 69:19]
  reg [31:0] writeMasterReg_Addr; // @[WriteNoBuffer.scala 72:27]
  reg [31:0] writeMasterReg_Data; // @[WriteNoBuffer.scala 72:27]
  reg [3:0] writeMasterReg_ByteEn; // @[WriteNoBuffer.scala 72:27]
  wire [1:0] wrPos = writeMasterReg_Addr[3:2]; // @[WriteNoBuffer.scala 82:34]
  wire [27:0] hi = writeMasterReg_Addr[31:4]; // @[WriteNoBuffer.scala 89:49]
  wire [31:0] _T_2 = {hi,4'h0}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_0 = cntReg == 2'h0 ? 3'h1 : io_readMaster_M_Cmd; // @[WriteNoBuffer.scala 87:30 WriteNoBuffer.scala 88:22 WriteNoBuffer.scala 80:14]
  wire [31:0] _GEN_1 = cntReg == 2'h0 ? _T_2 : io_readMaster_M_Addr; // @[WriteNoBuffer.scala 87:30 WriteNoBuffer.scala 89:23 WriteNoBuffer.scala 80:14]
  wire [3:0] _GEN_2 = cntReg == wrPos ? writeMasterReg_ByteEn : 4'h0; // @[WriteNoBuffer.scala 95:28 WriteNoBuffer.scala 96:29 WriteNoBuffer.scala 94:27]
  wire [1:0] _T_6 = cntReg + 2'h1; // @[WriteNoBuffer.scala 99:24]
  wire [1:0] _GEN_4 = cntReg == 2'h3 ? 2'h2 : state; // @[WriteNoBuffer.scala 101:44 WriteNoBuffer.scala 102:13 WriteNoBuffer.scala 68:18]
  wire [1:0] _GEN_5 = state == 2'h1 ? 2'h0 : io_slave_S_Resp; // @[WriteNoBuffer.scala 85:25 WriteNoBuffer.scala 86:26 WriteNoBuffer.scala 75:19]
  wire [1:0] _GEN_12 = state == 2'h1 ? _GEN_4 : state; // @[WriteNoBuffer.scala 85:25 WriteNoBuffer.scala 68:18]
  assign io_readMaster_S_Resp = state == 2'h2 ? 2'h0 : _GEN_5; // @[WriteNoBuffer.scala 105:29 WriteNoBuffer.scala 106:26]
  assign io_readMaster_S_Data = io_slave_S_Data; // @[WriteNoBuffer.scala 75:19]
  assign io_readMaster_S_CmdAccept = io_slave_S_CmdAccept; // @[WriteNoBuffer.scala 75:19]
  assign io_readMaster_S_DataAccept = io_slave_S_DataAccept; // @[WriteNoBuffer.scala 75:19]
  assign io_writeMaster_S_Resp = state == 2'h2 ? io_slave_S_Resp : 2'h0; // @[WriteNoBuffer.scala 105:29 WriteNoBuffer.scala 107:27 WriteNoBuffer.scala 77:25]
  assign io_slave_M_Cmd = state == 2'h1 ? _GEN_0 : io_readMaster_M_Cmd; // @[WriteNoBuffer.scala 85:25 WriteNoBuffer.scala 80:14]
  assign io_slave_M_Addr = state == 2'h1 ? _GEN_1 : io_readMaster_M_Addr; // @[WriteNoBuffer.scala 85:25 WriteNoBuffer.scala 80:14]
  assign io_slave_M_Data = state == 2'h1 ? writeMasterReg_Data : io_readMaster_M_Data; // @[WriteNoBuffer.scala 85:25 WriteNoBuffer.scala 93:21 WriteNoBuffer.scala 80:14]
  assign io_slave_M_DataValid = state == 2'h1 | io_readMaster_M_DataValid; // @[WriteNoBuffer.scala 85:25 WriteNoBuffer.scala 92:26 WriteNoBuffer.scala 80:14]
  assign io_slave_M_DataByteEn = state == 2'h1 ? _GEN_2 : io_readMaster_M_DataByteEn; // @[WriteNoBuffer.scala 85:25 WriteNoBuffer.scala 80:14]
  always @(posedge clock) begin
    if (reset) begin // @[WriteNoBuffer.scala 68:18]
      state <= 2'h0; // @[WriteNoBuffer.scala 68:18]
    end else if (io_writeMaster_M_Cmd == 3'h1) begin // @[WriteNoBuffer.scala 117:44]
      state <= 2'h1; // @[WriteNoBuffer.scala 118:11]
    end else if (state == 2'h2) begin // @[WriteNoBuffer.scala 105:29]
      if (io_slave_S_Resp != 2'h0) begin // @[WriteNoBuffer.scala 108:44]
        state <= 2'h0; // @[WriteNoBuffer.scala 109:13]
      end else begin
        state <= _GEN_12;
      end
    end else begin
      state <= _GEN_12;
    end
    if (reset) begin // @[WriteNoBuffer.scala 69:19]
      cntReg <= 2'h0; // @[WriteNoBuffer.scala 69:19]
    end else if (state == 2'h1) begin // @[WriteNoBuffer.scala 85:25]
      if (io_slave_S_DataAccept) begin // @[WriteNoBuffer.scala 98:45]
        cntReg <= _T_6; // @[WriteNoBuffer.scala 99:14]
      end
    end
    if (state != 2'h1) begin // @[WriteNoBuffer.scala 112:25]
      writeMasterReg_Addr <= io_writeMaster_M_Addr; // @[WriteNoBuffer.scala 113:20]
    end
    if (state != 2'h1) begin // @[WriteNoBuffer.scala 112:25]
      writeMasterReg_Data <= io_writeMaster_M_Data; // @[WriteNoBuffer.scala 113:20]
    end
    if (state != 2'h1) begin // @[WriteNoBuffer.scala 112:25]
      writeMasterReg_ByteEn <= io_writeMaster_M_ByteEn; // @[WriteNoBuffer.scala 113:20]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cntReg = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  writeMasterReg_Addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  writeMasterReg_Data = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  writeMasterReg_ByteEn = _RAND_4[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DataCache(
  input         clock,
  input         reset,
  input  [2:0]  io_master_M_Cmd,
  input  [31:0] io_master_M_Addr,
  input  [31:0] io_master_M_Data,
  input  [3:0]  io_master_M_ByteEn,
  input  [1:0]  io_master_M_AddrSpace,
  output [1:0]  io_master_S_Resp,
  output [31:0] io_master_S_Data,
  output [2:0]  io_slave_M_Cmd,
  output [31:0] io_slave_M_Addr,
  output [31:0] io_slave_M_Data,
  output        io_slave_M_DataValid,
  output [3:0]  io_slave_M_DataByteEn,
  input  [1:0]  io_slave_S_Resp,
  input  [31:0] io_slave_S_Data,
  input         io_slave_S_CmdAccept,
  input         io_slave_S_DataAccept,
  input         io_scIO_ena_in,
  input  [2:0]  io_scIO_exsc_op,
  input  [31:0] io_scIO_exsc_opData,
  input  [31:0] io_scIO_exsc_opOff,
  output [31:0] io_scIO_scex_stackTop,
  output [31:0] io_scIO_scex_memTop,
  output        io_scIO_illMem,
  output        io_scIO_stall,
  input         io_invalDCache
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  dm_clock; // @[DataCache.scala 44:13]
  wire  dm_reset; // @[DataCache.scala 44:13]
  wire [2:0] dm_io_master_M_Cmd; // @[DataCache.scala 44:13]
  wire [31:0] dm_io_master_M_Addr; // @[DataCache.scala 44:13]
  wire [31:0] dm_io_master_M_Data; // @[DataCache.scala 44:13]
  wire [3:0] dm_io_master_M_ByteEn; // @[DataCache.scala 44:13]
  wire [1:0] dm_io_master_S_Resp; // @[DataCache.scala 44:13]
  wire [31:0] dm_io_master_S_Data; // @[DataCache.scala 44:13]
  wire [2:0] dm_io_slave_M_Cmd; // @[DataCache.scala 44:13]
  wire [31:0] dm_io_slave_M_Addr; // @[DataCache.scala 44:13]
  wire [1:0] dm_io_slave_S_Resp; // @[DataCache.scala 44:13]
  wire [31:0] dm_io_slave_S_Data; // @[DataCache.scala 44:13]
  wire  dm_io_slave_S_CmdAccept; // @[DataCache.scala 44:13]
  wire  dm_io_invalidate; // @[DataCache.scala 44:13]
  wire  sc_clock; // @[DataCache.scala 66:18]
  wire  sc_reset; // @[DataCache.scala 66:18]
  wire  sc_io_ena_in; // @[DataCache.scala 66:18]
  wire [2:0] sc_io_exsc_op; // @[DataCache.scala 66:18]
  wire [31:0] sc_io_exsc_opData; // @[DataCache.scala 66:18]
  wire [31:0] sc_io_exsc_opOff; // @[DataCache.scala 66:18]
  wire [31:0] sc_io_scex_stackTop; // @[DataCache.scala 66:18]
  wire [31:0] sc_io_scex_memTop; // @[DataCache.scala 66:18]
  wire  sc_io_illMem; // @[DataCache.scala 66:18]
  wire  sc_io_stall; // @[DataCache.scala 66:18]
  wire [2:0] sc_io_fromCPU_M_Cmd; // @[DataCache.scala 66:18]
  wire [31:0] sc_io_fromCPU_M_Addr; // @[DataCache.scala 66:18]
  wire [31:0] sc_io_fromCPU_M_Data; // @[DataCache.scala 66:18]
  wire [3:0] sc_io_fromCPU_M_ByteEn; // @[DataCache.scala 66:18]
  wire [1:0] sc_io_fromCPU_S_Resp; // @[DataCache.scala 66:18]
  wire [31:0] sc_io_fromCPU_S_Data; // @[DataCache.scala 66:18]
  wire [2:0] sc_io_toMemory_M_Cmd; // @[DataCache.scala 66:18]
  wire [31:0] sc_io_toMemory_M_Addr; // @[DataCache.scala 66:18]
  wire [31:0] sc_io_toMemory_M_Data; // @[DataCache.scala 66:18]
  wire  sc_io_toMemory_M_DataValid; // @[DataCache.scala 66:18]
  wire [3:0] sc_io_toMemory_M_DataByteEn; // @[DataCache.scala 66:18]
  wire [1:0] sc_io_toMemory_S_Resp; // @[DataCache.scala 66:18]
  wire [31:0] sc_io_toMemory_S_Data; // @[DataCache.scala 66:18]
  wire  sc_io_toMemory_S_CmdAccept; // @[DataCache.scala 66:18]
  wire  bp_clock; // @[DataCache.scala 75:18]
  wire  bp_reset; // @[DataCache.scala 75:18]
  wire [2:0] bp_io_master_M_Cmd; // @[DataCache.scala 75:18]
  wire [31:0] bp_io_master_M_Addr; // @[DataCache.scala 75:18]
  wire [1:0] bp_io_master_S_Resp; // @[DataCache.scala 75:18]
  wire [31:0] bp_io_master_S_Data; // @[DataCache.scala 75:18]
  wire [2:0] bp_io_slave_M_Cmd; // @[DataCache.scala 75:18]
  wire [31:0] bp_io_slave_M_Addr; // @[DataCache.scala 75:18]
  wire [1:0] bp_io_slave_S_Resp; // @[DataCache.scala 75:18]
  wire [31:0] bp_io_slave_S_Data; // @[DataCache.scala 75:18]
  wire  bp_io_slave_S_CmdAccept; // @[DataCache.scala 75:18]
  wire [2:0] burstReadBus1_io_master_M_Cmd; // @[DataCache.scala 81:29]
  wire [31:0] burstReadBus1_io_master_M_Addr; // @[DataCache.scala 81:29]
  wire [31:0] burstReadBus1_io_master_M_Data; // @[DataCache.scala 81:29]
  wire  burstReadBus1_io_master_M_DataValid; // @[DataCache.scala 81:29]
  wire [3:0] burstReadBus1_io_master_M_DataByteEn; // @[DataCache.scala 81:29]
  wire [1:0] burstReadBus1_io_master_S_Resp; // @[DataCache.scala 81:29]
  wire [31:0] burstReadBus1_io_master_S_Data; // @[DataCache.scala 81:29]
  wire  burstReadBus1_io_master_S_CmdAccept; // @[DataCache.scala 81:29]
  wire  burstReadBus1_io_master_S_DataAccept; // @[DataCache.scala 81:29]
  wire [2:0] burstReadBus1_io_slave_M_Cmd; // @[DataCache.scala 81:29]
  wire [31:0] burstReadBus1_io_slave_M_Addr; // @[DataCache.scala 81:29]
  wire [31:0] burstReadBus1_io_slave_M_Data; // @[DataCache.scala 81:29]
  wire  burstReadBus1_io_slave_M_DataValid; // @[DataCache.scala 81:29]
  wire [3:0] burstReadBus1_io_slave_M_DataByteEn; // @[DataCache.scala 81:29]
  wire [1:0] burstReadBus1_io_slave_S_Resp; // @[DataCache.scala 81:29]
  wire [31:0] burstReadBus1_io_slave_S_Data; // @[DataCache.scala 81:29]
  wire  burstReadBus1_io_slave_S_CmdAccept; // @[DataCache.scala 81:29]
  wire  burstReadBus1_io_slave_S_DataAccept; // @[DataCache.scala 81:29]
  wire [2:0] burstReadBus2_io_master_M_Cmd; // @[DataCache.scala 84:29]
  wire [31:0] burstReadBus2_io_master_M_Addr; // @[DataCache.scala 84:29]
  wire [31:0] burstReadBus2_io_master_M_Data; // @[DataCache.scala 84:29]
  wire  burstReadBus2_io_master_M_DataValid; // @[DataCache.scala 84:29]
  wire [3:0] burstReadBus2_io_master_M_DataByteEn; // @[DataCache.scala 84:29]
  wire [1:0] burstReadBus2_io_master_S_Resp; // @[DataCache.scala 84:29]
  wire [31:0] burstReadBus2_io_master_S_Data; // @[DataCache.scala 84:29]
  wire  burstReadBus2_io_master_S_CmdAccept; // @[DataCache.scala 84:29]
  wire  burstReadBus2_io_master_S_DataAccept; // @[DataCache.scala 84:29]
  wire [2:0] burstReadBus2_io_slave_M_Cmd; // @[DataCache.scala 84:29]
  wire [31:0] burstReadBus2_io_slave_M_Addr; // @[DataCache.scala 84:29]
  wire [31:0] burstReadBus2_io_slave_M_Data; // @[DataCache.scala 84:29]
  wire  burstReadBus2_io_slave_M_DataValid; // @[DataCache.scala 84:29]
  wire [3:0] burstReadBus2_io_slave_M_DataByteEn; // @[DataCache.scala 84:29]
  wire [1:0] burstReadBus2_io_slave_S_Resp; // @[DataCache.scala 84:29]
  wire [31:0] burstReadBus2_io_slave_S_Data; // @[DataCache.scala 84:29]
  wire  burstReadBus2_io_slave_S_CmdAccept; // @[DataCache.scala 84:29]
  wire  burstReadBus2_io_slave_S_DataAccept; // @[DataCache.scala 84:29]
  wire  wc_clock; // @[DataCache.scala 88:18]
  wire  wc_reset; // @[DataCache.scala 88:18]
  wire [2:0] wc_io_readMaster_M_Cmd; // @[DataCache.scala 88:18]
  wire [31:0] wc_io_readMaster_M_Addr; // @[DataCache.scala 88:18]
  wire [31:0] wc_io_readMaster_M_Data; // @[DataCache.scala 88:18]
  wire  wc_io_readMaster_M_DataValid; // @[DataCache.scala 88:18]
  wire [3:0] wc_io_readMaster_M_DataByteEn; // @[DataCache.scala 88:18]
  wire [1:0] wc_io_readMaster_S_Resp; // @[DataCache.scala 88:18]
  wire [31:0] wc_io_readMaster_S_Data; // @[DataCache.scala 88:18]
  wire  wc_io_readMaster_S_CmdAccept; // @[DataCache.scala 88:18]
  wire  wc_io_readMaster_S_DataAccept; // @[DataCache.scala 88:18]
  wire [2:0] wc_io_writeMaster_M_Cmd; // @[DataCache.scala 88:18]
  wire [31:0] wc_io_writeMaster_M_Addr; // @[DataCache.scala 88:18]
  wire [31:0] wc_io_writeMaster_M_Data; // @[DataCache.scala 88:18]
  wire [3:0] wc_io_writeMaster_M_ByteEn; // @[DataCache.scala 88:18]
  wire [1:0] wc_io_writeMaster_S_Resp; // @[DataCache.scala 88:18]
  wire [2:0] wc_io_slave_M_Cmd; // @[DataCache.scala 88:18]
  wire [31:0] wc_io_slave_M_Addr; // @[DataCache.scala 88:18]
  wire [31:0] wc_io_slave_M_Data; // @[DataCache.scala 88:18]
  wire  wc_io_slave_M_DataValid; // @[DataCache.scala 88:18]
  wire [3:0] wc_io_slave_M_DataByteEn; // @[DataCache.scala 88:18]
  wire [1:0] wc_io_slave_S_Resp; // @[DataCache.scala 88:18]
  wire [31:0] wc_io_slave_S_Data; // @[DataCache.scala 88:18]
  wire  wc_io_slave_S_CmdAccept; // @[DataCache.scala 88:18]
  wire  wc_io_slave_S_DataAccept; // @[DataCache.scala 88:18]
  wire  selDC = io_master_M_AddrSpace == 2'h2; // @[DataCache.scala 30:62]
  reg  selDCReg; // @[DataCache.scala 31:21]
  wire  selSC = io_master_M_AddrSpace == 2'h0; // @[DataCache.scala 32:37]
  reg  selSCReg; // @[DataCache.scala 33:21]
  wire  _T_3 = io_master_M_Cmd == 3'h1; // @[DataCache.scala 60:46]
  wire  _T_9 = ~selSC; // @[DataCache.scala 77:39]
  reg  REG; // @[OcpBurst.scala 144:24]
  wire  _T_14 = bp_io_slave_M_Cmd != 3'h0 | REG; // @[OcpBurst.scala 147:25]
  wire  _T_15 = dm_io_slave_M_Cmd != 3'h0 ? 1'h0 : _T_14; // @[OcpBurst.scala 146:18]
  reg  REG_1; // @[OcpBurst.scala 144:24]
  wire  _T_20 = burstReadBus1_io_master_M_Cmd != 3'h0 | REG_1; // @[OcpBurst.scala 147:25]
  wire  _T_21 = sc_io_toMemory_M_Cmd != 3'h0 ? 1'h0 : _T_20; // @[OcpBurst.scala 146:18]
  wire [31:0] _GEN_16 = selDCReg ? dm_io_master_S_Data : bp_io_master_S_Data; // @[DataCache.scala 99:18 DataCache.scala 99:37 DataCache.scala 98:20]
  wire [1:0] _T_29 = dm_io_master_S_Resp | sc_io_fromCPU_S_Resp; // @[DataCache.scala 103:32]
  wire [1:0] _T_30 = _T_29 | bp_io_master_S_Resp; // @[DataCache.scala 103:43]
  DirectMappedCache dm ( // @[DataCache.scala 44:13]
    .clock(dm_clock),
    .reset(dm_reset),
    .io_master_M_Cmd(dm_io_master_M_Cmd),
    .io_master_M_Addr(dm_io_master_M_Addr),
    .io_master_M_Data(dm_io_master_M_Data),
    .io_master_M_ByteEn(dm_io_master_M_ByteEn),
    .io_master_S_Resp(dm_io_master_S_Resp),
    .io_master_S_Data(dm_io_master_S_Data),
    .io_slave_M_Cmd(dm_io_slave_M_Cmd),
    .io_slave_M_Addr(dm_io_slave_M_Addr),
    .io_slave_S_Resp(dm_io_slave_S_Resp),
    .io_slave_S_Data(dm_io_slave_S_Data),
    .io_slave_S_CmdAccept(dm_io_slave_S_CmdAccept),
    .io_invalidate(dm_io_invalidate)
  );
  StackCache sc ( // @[DataCache.scala 66:18]
    .clock(sc_clock),
    .reset(sc_reset),
    .io_ena_in(sc_io_ena_in),
    .io_exsc_op(sc_io_exsc_op),
    .io_exsc_opData(sc_io_exsc_opData),
    .io_exsc_opOff(sc_io_exsc_opOff),
    .io_scex_stackTop(sc_io_scex_stackTop),
    .io_scex_memTop(sc_io_scex_memTop),
    .io_illMem(sc_io_illMem),
    .io_stall(sc_io_stall),
    .io_fromCPU_M_Cmd(sc_io_fromCPU_M_Cmd),
    .io_fromCPU_M_Addr(sc_io_fromCPU_M_Addr),
    .io_fromCPU_M_Data(sc_io_fromCPU_M_Data),
    .io_fromCPU_M_ByteEn(sc_io_fromCPU_M_ByteEn),
    .io_fromCPU_S_Resp(sc_io_fromCPU_S_Resp),
    .io_fromCPU_S_Data(sc_io_fromCPU_S_Data),
    .io_toMemory_M_Cmd(sc_io_toMemory_M_Cmd),
    .io_toMemory_M_Addr(sc_io_toMemory_M_Addr),
    .io_toMemory_M_Data(sc_io_toMemory_M_Data),
    .io_toMemory_M_DataValid(sc_io_toMemory_M_DataValid),
    .io_toMemory_M_DataByteEn(sc_io_toMemory_M_DataByteEn),
    .io_toMemory_S_Resp(sc_io_toMemory_S_Resp),
    .io_toMemory_S_Data(sc_io_toMemory_S_Data),
    .io_toMemory_S_CmdAccept(sc_io_toMemory_S_CmdAccept)
  );
  NullCache bp ( // @[DataCache.scala 75:18]
    .clock(bp_clock),
    .reset(bp_reset),
    .io_master_M_Cmd(bp_io_master_M_Cmd),
    .io_master_M_Addr(bp_io_master_M_Addr),
    .io_master_S_Resp(bp_io_master_S_Resp),
    .io_master_S_Data(bp_io_master_S_Data),
    .io_slave_M_Cmd(bp_io_slave_M_Cmd),
    .io_slave_M_Addr(bp_io_slave_M_Addr),
    .io_slave_S_Resp(bp_io_slave_S_Resp),
    .io_slave_S_Data(bp_io_slave_S_Data),
    .io_slave_S_CmdAccept(bp_io_slave_S_CmdAccept)
  );
  OcpBurstBus burstReadBus1 ( // @[DataCache.scala 81:29]
    .io_master_M_Cmd(burstReadBus1_io_master_M_Cmd),
    .io_master_M_Addr(burstReadBus1_io_master_M_Addr),
    .io_master_M_Data(burstReadBus1_io_master_M_Data),
    .io_master_M_DataValid(burstReadBus1_io_master_M_DataValid),
    .io_master_M_DataByteEn(burstReadBus1_io_master_M_DataByteEn),
    .io_master_S_Resp(burstReadBus1_io_master_S_Resp),
    .io_master_S_Data(burstReadBus1_io_master_S_Data),
    .io_master_S_CmdAccept(burstReadBus1_io_master_S_CmdAccept),
    .io_master_S_DataAccept(burstReadBus1_io_master_S_DataAccept),
    .io_slave_M_Cmd(burstReadBus1_io_slave_M_Cmd),
    .io_slave_M_Addr(burstReadBus1_io_slave_M_Addr),
    .io_slave_M_Data(burstReadBus1_io_slave_M_Data),
    .io_slave_M_DataValid(burstReadBus1_io_slave_M_DataValid),
    .io_slave_M_DataByteEn(burstReadBus1_io_slave_M_DataByteEn),
    .io_slave_S_Resp(burstReadBus1_io_slave_S_Resp),
    .io_slave_S_Data(burstReadBus1_io_slave_S_Data),
    .io_slave_S_CmdAccept(burstReadBus1_io_slave_S_CmdAccept),
    .io_slave_S_DataAccept(burstReadBus1_io_slave_S_DataAccept)
  );
  OcpBurstBus burstReadBus2 ( // @[DataCache.scala 84:29]
    .io_master_M_Cmd(burstReadBus2_io_master_M_Cmd),
    .io_master_M_Addr(burstReadBus2_io_master_M_Addr),
    .io_master_M_Data(burstReadBus2_io_master_M_Data),
    .io_master_M_DataValid(burstReadBus2_io_master_M_DataValid),
    .io_master_M_DataByteEn(burstReadBus2_io_master_M_DataByteEn),
    .io_master_S_Resp(burstReadBus2_io_master_S_Resp),
    .io_master_S_Data(burstReadBus2_io_master_S_Data),
    .io_master_S_CmdAccept(burstReadBus2_io_master_S_CmdAccept),
    .io_master_S_DataAccept(burstReadBus2_io_master_S_DataAccept),
    .io_slave_M_Cmd(burstReadBus2_io_slave_M_Cmd),
    .io_slave_M_Addr(burstReadBus2_io_slave_M_Addr),
    .io_slave_M_Data(burstReadBus2_io_slave_M_Data),
    .io_slave_M_DataValid(burstReadBus2_io_slave_M_DataValid),
    .io_slave_M_DataByteEn(burstReadBus2_io_slave_M_DataByteEn),
    .io_slave_S_Resp(burstReadBus2_io_slave_S_Resp),
    .io_slave_S_Data(burstReadBus2_io_slave_S_Data),
    .io_slave_S_CmdAccept(burstReadBus2_io_slave_S_CmdAccept),
    .io_slave_S_DataAccept(burstReadBus2_io_slave_S_DataAccept)
  );
  WriteNoBuffer wc ( // @[DataCache.scala 88:18]
    .clock(wc_clock),
    .reset(wc_reset),
    .io_readMaster_M_Cmd(wc_io_readMaster_M_Cmd),
    .io_readMaster_M_Addr(wc_io_readMaster_M_Addr),
    .io_readMaster_M_Data(wc_io_readMaster_M_Data),
    .io_readMaster_M_DataValid(wc_io_readMaster_M_DataValid),
    .io_readMaster_M_DataByteEn(wc_io_readMaster_M_DataByteEn),
    .io_readMaster_S_Resp(wc_io_readMaster_S_Resp),
    .io_readMaster_S_Data(wc_io_readMaster_S_Data),
    .io_readMaster_S_CmdAccept(wc_io_readMaster_S_CmdAccept),
    .io_readMaster_S_DataAccept(wc_io_readMaster_S_DataAccept),
    .io_writeMaster_M_Cmd(wc_io_writeMaster_M_Cmd),
    .io_writeMaster_M_Addr(wc_io_writeMaster_M_Addr),
    .io_writeMaster_M_Data(wc_io_writeMaster_M_Data),
    .io_writeMaster_M_ByteEn(wc_io_writeMaster_M_ByteEn),
    .io_writeMaster_S_Resp(wc_io_writeMaster_S_Resp),
    .io_slave_M_Cmd(wc_io_slave_M_Cmd),
    .io_slave_M_Addr(wc_io_slave_M_Addr),
    .io_slave_M_Data(wc_io_slave_M_Data),
    .io_slave_M_DataValid(wc_io_slave_M_DataValid),
    .io_slave_M_DataByteEn(wc_io_slave_M_DataByteEn),
    .io_slave_S_Resp(wc_io_slave_S_Resp),
    .io_slave_S_Data(wc_io_slave_S_Data),
    .io_slave_S_CmdAccept(wc_io_slave_S_CmdAccept),
    .io_slave_S_DataAccept(wc_io_slave_S_DataAccept)
  );
  assign io_master_S_Resp = _T_30 | wc_io_writeMaster_S_Resp; // @[DataCache.scala 103:54]
  assign io_master_S_Data = selSCReg ? sc_io_fromCPU_S_Data : _GEN_16; // @[DataCache.scala 100:18 DataCache.scala 100:37]
  assign io_slave_M_Cmd = wc_io_slave_M_Cmd; // @[DataCache.scala 95:12]
  assign io_slave_M_Addr = wc_io_slave_M_Addr; // @[DataCache.scala 95:12]
  assign io_slave_M_Data = wc_io_slave_M_Data; // @[DataCache.scala 95:12]
  assign io_slave_M_DataValid = wc_io_slave_M_DataValid; // @[DataCache.scala 95:12]
  assign io_slave_M_DataByteEn = wc_io_slave_M_DataByteEn; // @[DataCache.scala 95:12]
  assign io_scIO_scex_stackTop = sc_io_scex_stackTop; // @[DataCache.scala 67:11]
  assign io_scIO_scex_memTop = sc_io_scex_memTop; // @[DataCache.scala 67:11]
  assign io_scIO_illMem = sc_io_illMem; // @[DataCache.scala 67:11]
  assign io_scIO_stall = sc_io_stall; // @[DataCache.scala 67:11]
  assign dm_clock = clock;
  assign dm_reset = reset;
  assign dm_io_master_M_Cmd = selDC | _T_3 ? io_master_M_Cmd : 3'h0; // @[DataCache.scala 58:28]
  assign dm_io_master_M_Addr = io_master_M_Addr; // @[DataCache.scala 57:18]
  assign dm_io_master_M_Data = io_master_M_Data; // @[DataCache.scala 57:18]
  assign dm_io_master_M_ByteEn = io_master_M_ByteEn; // @[DataCache.scala 57:18]
  assign dm_io_slave_S_Resp = REG ? 2'h0 : burstReadBus1_io_slave_S_Resp; // @[OcpBurst.scala 159:21 OcpBurst.scala 160:17 OcpBurst.scala 157:10]
  assign dm_io_slave_S_Data = burstReadBus1_io_slave_S_Data; // @[OcpBurst.scala 157:10]
  assign dm_io_slave_S_CmdAccept = burstReadBus1_io_slave_S_CmdAccept; // @[OcpBurst.scala 157:10]
  assign dm_io_invalidate = io_invalDCache; // @[DataCache.scala 62:20]
  assign sc_clock = clock;
  assign sc_reset = reset;
  assign sc_io_ena_in = io_scIO_ena_in; // @[DataCache.scala 67:11]
  assign sc_io_exsc_op = io_scIO_exsc_op; // @[DataCache.scala 67:11]
  assign sc_io_exsc_opData = io_scIO_exsc_opData; // @[DataCache.scala 67:11]
  assign sc_io_exsc_opOff = io_scIO_exsc_opOff; // @[DataCache.scala 67:11]
  assign sc_io_fromCPU_M_Cmd = selSC ? io_master_M_Cmd : 3'h0; // @[DataCache.scala 71:29]
  assign sc_io_fromCPU_M_Addr = io_master_M_Addr; // @[DataCache.scala 70:19]
  assign sc_io_fromCPU_M_Data = io_master_M_Data; // @[DataCache.scala 70:19]
  assign sc_io_fromCPU_M_ByteEn = io_master_M_ByteEn; // @[DataCache.scala 70:19]
  assign sc_io_toMemory_S_Resp = REG_1 ? 2'h0 : burstReadBus2_io_slave_S_Resp; // @[OcpBurst.scala 159:21 OcpBurst.scala 160:17 OcpBurst.scala 157:10]
  assign sc_io_toMemory_S_Data = burstReadBus2_io_slave_S_Data; // @[OcpBurst.scala 157:10]
  assign sc_io_toMemory_S_CmdAccept = burstReadBus2_io_slave_S_CmdAccept; // @[OcpBurst.scala 157:10]
  assign bp_clock = clock;
  assign bp_reset = reset;
  assign bp_io_master_M_Cmd = ~selDC & ~selSC ? io_master_M_Cmd : 3'h0; // @[DataCache.scala 77:28]
  assign bp_io_master_M_Addr = io_master_M_Addr; // @[DataCache.scala 76:18]
  assign bp_io_slave_S_Resp = REG ? burstReadBus1_io_slave_S_Resp : 2'h0; // @[OcpBurst.scala 159:21 OcpBurst.scala 156:11 OcpBurst.scala 163:18]
  assign bp_io_slave_S_Data = burstReadBus1_io_slave_S_Data; // @[OcpBurst.scala 156:11]
  assign bp_io_slave_S_CmdAccept = burstReadBus1_io_slave_S_CmdAccept; // @[OcpBurst.scala 156:11]
  assign burstReadBus1_io_master_S_Resp = REG_1 ? burstReadBus2_io_slave_S_Resp : 2'h0; // @[OcpBurst.scala 159:21 OcpBurst.scala 156:11 OcpBurst.scala 163:18]
  assign burstReadBus1_io_master_S_Data = burstReadBus2_io_slave_S_Data; // @[OcpBurst.scala 156:11]
  assign burstReadBus1_io_master_S_CmdAccept = burstReadBus2_io_slave_S_CmdAccept; // @[OcpBurst.scala 156:11]
  assign burstReadBus1_io_master_S_DataAccept = burstReadBus2_io_slave_S_DataAccept; // @[OcpBurst.scala 156:11]
  assign burstReadBus1_io_slave_M_Cmd = bp_io_slave_M_Cmd | dm_io_slave_M_Cmd; // @[OcpBurst.scala 154:31]
  assign burstReadBus1_io_slave_M_Addr = _T_15 ? bp_io_slave_M_Addr : dm_io_slave_M_Addr; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign burstReadBus1_io_slave_M_Data = 32'h0; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign burstReadBus1_io_slave_M_DataValid = 1'h0; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign burstReadBus1_io_slave_M_DataByteEn = 4'h0; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign burstReadBus2_io_master_S_Resp = wc_io_readMaster_S_Resp; // @[DataCache.scala 90:29]
  assign burstReadBus2_io_master_S_Data = wc_io_readMaster_S_Data; // @[DataCache.scala 90:29]
  assign burstReadBus2_io_master_S_CmdAccept = wc_io_readMaster_S_CmdAccept; // @[DataCache.scala 90:29]
  assign burstReadBus2_io_master_S_DataAccept = wc_io_readMaster_S_DataAccept; // @[DataCache.scala 90:29]
  assign burstReadBus2_io_slave_M_Cmd = burstReadBus1_io_master_M_Cmd | sc_io_toMemory_M_Cmd; // @[OcpBurst.scala 154:31]
  assign burstReadBus2_io_slave_M_Addr = _T_21 ? burstReadBus1_io_master_M_Addr : sc_io_toMemory_M_Addr; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign burstReadBus2_io_slave_M_Data = _T_21 ? burstReadBus1_io_master_M_Data : sc_io_toMemory_M_Data; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign burstReadBus2_io_slave_M_DataValid = _T_21 ? burstReadBus1_io_master_M_DataValid : sc_io_toMemory_M_DataValid; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign burstReadBus2_io_slave_M_DataByteEn = _T_21 ? burstReadBus1_io_master_M_DataByteEn :
    sc_io_toMemory_M_DataByteEn; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign wc_clock = clock;
  assign wc_reset = reset;
  assign wc_io_readMaster_M_Cmd = burstReadBus2_io_master_M_Cmd; // @[DataCache.scala 89:22]
  assign wc_io_readMaster_M_Addr = burstReadBus2_io_master_M_Addr; // @[DataCache.scala 89:22]
  assign wc_io_readMaster_M_Data = burstReadBus2_io_master_M_Data; // @[DataCache.scala 89:22]
  assign wc_io_readMaster_M_DataValid = burstReadBus2_io_master_M_DataValid; // @[DataCache.scala 89:22]
  assign wc_io_readMaster_M_DataByteEn = burstReadBus2_io_master_M_DataByteEn; // @[DataCache.scala 89:22]
  assign wc_io_writeMaster_M_Cmd = _T_9 ? io_master_M_Cmd : 3'h0; // @[DataCache.scala 92:33]
  assign wc_io_writeMaster_M_Addr = io_master_M_Addr; // @[DataCache.scala 91:23]
  assign wc_io_writeMaster_M_Data = io_master_M_Data; // @[DataCache.scala 91:23]
  assign wc_io_writeMaster_M_ByteEn = io_master_M_ByteEn; // @[DataCache.scala 91:23]
  assign wc_io_slave_S_Resp = io_slave_S_Resp; // @[DataCache.scala 95:12]
  assign wc_io_slave_S_Data = io_slave_S_Data; // @[DataCache.scala 95:12]
  assign wc_io_slave_S_CmdAccept = io_slave_S_CmdAccept; // @[DataCache.scala 95:12]
  assign wc_io_slave_S_DataAccept = io_slave_S_DataAccept; // @[DataCache.scala 95:12]
  always @(posedge clock) begin
    if (io_master_M_Cmd != 3'h0) begin // @[DataCache.scala 34:41]
      selDCReg <= selDC; // @[DataCache.scala 35:14]
    end
    if (io_master_M_Cmd != 3'h0) begin // @[DataCache.scala 34:41]
      selSCReg <= selSC; // @[DataCache.scala 36:14]
    end
    if (dm_io_slave_M_Cmd != 3'h0) begin // @[OcpBurst.scala 146:18]
      REG <= 1'h0;
    end else begin
      REG <= _T_14;
    end
    if (sc_io_toMemory_M_Cmd != 3'h0) begin // @[OcpBurst.scala 146:18]
      REG_1 <= 1'h0;
    end else begin
      REG_1 <= _T_20;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  selDCReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  selSCReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_1 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module NoMemoryManagement(
  input  [2:0]  io_virt_M_Cmd,
  input  [31:0] io_virt_M_Addr,
  input  [31:0] io_virt_M_Data,
  input         io_virt_M_DataValid,
  input  [3:0]  io_virt_M_DataByteEn,
  output [1:0]  io_virt_S_Resp,
  output [31:0] io_virt_S_Data,
  output [2:0]  io_phys_M_Cmd,
  output [20:0] io_phys_M_Addr,
  output [31:0] io_phys_M_Data,
  output        io_phys_M_DataValid,
  output [3:0]  io_phys_M_DataByteEn,
  input  [1:0]  io_phys_S_Resp,
  input  [31:0] io_phys_S_Data
);
  assign io_virt_S_Resp = io_phys_S_Resp; // @[NoMemoryManagement.scala 17:13]
  assign io_virt_S_Data = io_phys_S_Data; // @[NoMemoryManagement.scala 17:13]
  assign io_phys_M_Cmd = io_virt_M_Cmd; // @[NoMemoryManagement.scala 16:13]
  assign io_phys_M_Addr = io_virt_M_Addr[20:0]; // @[NoMemoryManagement.scala 16:13]
  assign io_phys_M_Data = io_virt_M_Data; // @[NoMemoryManagement.scala 16:13]
  assign io_phys_M_DataValid = io_virt_M_DataValid; // @[NoMemoryManagement.scala 16:13]
  assign io_phys_M_DataByteEn = io_virt_M_DataByteEn; // @[NoMemoryManagement.scala 16:13]
endmodule
module PatmosCore(
  input         clock,
  input         reset,
  input         io_interrupts_0,
  input         io_interrupts_1,
  input         io_interrupts_2,
  input         io_interrupts_3,
  input         io_interrupts_4,
  input         io_interrupts_5,
  output [2:0]  io_memPort_M_Cmd,
  output [20:0] io_memPort_M_Addr,
  output [31:0] io_memPort_M_Data,
  output        io_memPort_M_DataValid,
  output [3:0]  io_memPort_M_DataByteEn,
  input  [1:0]  io_memPort_S_Resp,
  input  [31:0] io_memPort_S_Data,
  output [2:0]  io_memInOut_M_Cmd,
  output [31:0] io_memInOut_M_Addr,
  output [31:0] io_memInOut_M_Data,
  output [3:0]  io_memInOut_M_ByteEn,
  input  [1:0]  io_memInOut_S_Resp,
  input  [31:0] io_memInOut_S_Data,
  input  [2:0]  io_excInOut_M_Cmd,
  input  [31:0] io_excInOut_M_Addr,
  input  [31:0] io_excInOut_M_Data,
  output [1:0]  io_excInOut_S_Resp,
  output [31:0] io_excInOut_S_Data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  icache_clock; // @[Patmos.scala 44:13]
  wire  icache_reset; // @[Patmos.scala 44:13]
  wire  icache_io_ena_out; // @[Patmos.scala 44:13]
  wire  icache_io_ena_in; // @[Patmos.scala 44:13]
  wire  icache_io_invalidate; // @[Patmos.scala 44:13]
  wire [31:0] icache_io_feicache_addrEven; // @[Patmos.scala 44:13]
  wire [31:0] icache_io_feicache_addrOdd; // @[Patmos.scala 44:13]
  wire  icache_io_exicache_doCallRet; // @[Patmos.scala 44:13]
  wire [31:0] icache_io_exicache_callRetBase; // @[Patmos.scala 44:13]
  wire [31:0] icache_io_exicache_callRetAddr; // @[Patmos.scala 44:13]
  wire [31:0] icache_io_icachefe_instrEven; // @[Patmos.scala 44:13]
  wire [31:0] icache_io_icachefe_instrOdd; // @[Patmos.scala 44:13]
  wire [31:0] icache_io_icachefe_base; // @[Patmos.scala 44:13]
  wire [10:0] icache_io_icachefe_relBase; // @[Patmos.scala 44:13]
  wire [11:0] icache_io_icachefe_relPc; // @[Patmos.scala 44:13]
  wire [31:0] icache_io_icachefe_reloc; // @[Patmos.scala 44:13]
  wire [1:0] icache_io_icachefe_memSel; // @[Patmos.scala 44:13]
  wire [2:0] icache_io_ocp_port_M_Cmd; // @[Patmos.scala 44:13]
  wire [31:0] icache_io_ocp_port_M_Addr; // @[Patmos.scala 44:13]
  wire [1:0] icache_io_ocp_port_S_Resp; // @[Patmos.scala 44:13]
  wire [31:0] icache_io_ocp_port_S_Data; // @[Patmos.scala 44:13]
  wire  icache_io_ocp_port_S_CmdAccept; // @[Patmos.scala 44:13]
  wire  icache_io_illMem; // @[Patmos.scala 44:13]
  wire  fetch_clock; // @[Patmos.scala 56:21]
  wire  fetch_reset; // @[Patmos.scala 56:21]
  wire  fetch_io_ena; // @[Patmos.scala 56:21]
  wire [31:0] fetch_io_fedec_instr_a; // @[Patmos.scala 56:21]
  wire [31:0] fetch_io_fedec_instr_b; // @[Patmos.scala 56:21]
  wire [29:0] fetch_io_fedec_pc; // @[Patmos.scala 56:21]
  wire [29:0] fetch_io_fedec_base; // @[Patmos.scala 56:21]
  wire [31:0] fetch_io_fedec_reloc; // @[Patmos.scala 56:21]
  wire [29:0] fetch_io_fedec_relPc; // @[Patmos.scala 56:21]
  wire [29:0] fetch_io_feex_pc; // @[Patmos.scala 56:21]
  wire  fetch_io_exfe_doBranch; // @[Patmos.scala 56:21]
  wire [29:0] fetch_io_exfe_branchPc; // @[Patmos.scala 56:21]
  wire  fetch_io_memfe_doCallRet; // @[Patmos.scala 56:21]
  wire  fetch_io_memfe_store; // @[Patmos.scala 56:21]
  wire [31:0] fetch_io_memfe_addr; // @[Patmos.scala 56:21]
  wire [31:0] fetch_io_memfe_data; // @[Patmos.scala 56:21]
  wire [31:0] fetch_io_feicache_addrEven; // @[Patmos.scala 56:21]
  wire [31:0] fetch_io_feicache_addrOdd; // @[Patmos.scala 56:21]
  wire [31:0] fetch_io_icachefe_instrEven; // @[Patmos.scala 56:21]
  wire [31:0] fetch_io_icachefe_instrOdd; // @[Patmos.scala 56:21]
  wire [31:0] fetch_io_icachefe_base; // @[Patmos.scala 56:21]
  wire [10:0] fetch_io_icachefe_relBase; // @[Patmos.scala 56:21]
  wire [11:0] fetch_io_icachefe_relPc; // @[Patmos.scala 56:21]
  wire [31:0] fetch_io_icachefe_reloc; // @[Patmos.scala 56:21]
  wire [1:0] fetch_io_icachefe_memSel; // @[Patmos.scala 56:21]
  wire  decode_clock; // @[Patmos.scala 57:22]
  wire  decode_reset; // @[Patmos.scala 57:22]
  wire  decode_io_ena; // @[Patmos.scala 57:22]
  wire  decode_io_flush; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_fedec_instr_a; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_fedec_instr_b; // @[Patmos.scala 57:22]
  wire [29:0] decode_io_fedec_pc; // @[Patmos.scala 57:22]
  wire [29:0] decode_io_fedec_base; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_fedec_reloc; // @[Patmos.scala 57:22]
  wire [29:0] decode_io_fedec_relPc; // @[Patmos.scala 57:22]
  wire [29:0] decode_io_decex_base; // @[Patmos.scala 57:22]
  wire [29:0] decode_io_decex_relPc; // @[Patmos.scala 57:22]
  wire [3:0] decode_io_decex_pred_0; // @[Patmos.scala 57:22]
  wire [3:0] decode_io_decex_pred_1; // @[Patmos.scala 57:22]
  wire [3:0] decode_io_decex_aluOp_0_func; // @[Patmos.scala 57:22]
  wire  decode_io_decex_aluOp_0_isMul; // @[Patmos.scala 57:22]
  wire  decode_io_decex_aluOp_0_isCmp; // @[Patmos.scala 57:22]
  wire  decode_io_decex_aluOp_0_isPred; // @[Patmos.scala 57:22]
  wire  decode_io_decex_aluOp_0_isBCpy; // @[Patmos.scala 57:22]
  wire  decode_io_decex_aluOp_0_isMTS; // @[Patmos.scala 57:22]
  wire  decode_io_decex_aluOp_0_isMFS; // @[Patmos.scala 57:22]
  wire [3:0] decode_io_decex_aluOp_1_func; // @[Patmos.scala 57:22]
  wire  decode_io_decex_aluOp_1_isCmp; // @[Patmos.scala 57:22]
  wire  decode_io_decex_aluOp_1_isPred; // @[Patmos.scala 57:22]
  wire  decode_io_decex_aluOp_1_isBCpy; // @[Patmos.scala 57:22]
  wire  decode_io_decex_aluOp_1_isMTS; // @[Patmos.scala 57:22]
  wire  decode_io_decex_aluOp_1_isMFS; // @[Patmos.scala 57:22]
  wire [1:0] decode_io_decex_predOp_0_func; // @[Patmos.scala 57:22]
  wire [2:0] decode_io_decex_predOp_0_dest; // @[Patmos.scala 57:22]
  wire [3:0] decode_io_decex_predOp_0_s1Addr; // @[Patmos.scala 57:22]
  wire [3:0] decode_io_decex_predOp_0_s2Addr; // @[Patmos.scala 57:22]
  wire [1:0] decode_io_decex_predOp_1_func; // @[Patmos.scala 57:22]
  wire [2:0] decode_io_decex_predOp_1_dest; // @[Patmos.scala 57:22]
  wire [3:0] decode_io_decex_predOp_1_s1Addr; // @[Patmos.scala 57:22]
  wire [3:0] decode_io_decex_predOp_1_s2Addr; // @[Patmos.scala 57:22]
  wire  decode_io_decex_jmpOp_branch; // @[Patmos.scala 57:22]
  wire [29:0] decode_io_decex_jmpOp_target; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_decex_jmpOp_reloc; // @[Patmos.scala 57:22]
  wire  decode_io_decex_memOp_load; // @[Patmos.scala 57:22]
  wire  decode_io_decex_memOp_store; // @[Patmos.scala 57:22]
  wire  decode_io_decex_memOp_hword; // @[Patmos.scala 57:22]
  wire  decode_io_decex_memOp_byte; // @[Patmos.scala 57:22]
  wire  decode_io_decex_memOp_zext; // @[Patmos.scala 57:22]
  wire [1:0] decode_io_decex_memOp_typ; // @[Patmos.scala 57:22]
  wire [2:0] decode_io_decex_stackOp; // @[Patmos.scala 57:22]
  wire [4:0] decode_io_decex_rsAddr_0; // @[Patmos.scala 57:22]
  wire [4:0] decode_io_decex_rsAddr_1; // @[Patmos.scala 57:22]
  wire [4:0] decode_io_decex_rsAddr_2; // @[Patmos.scala 57:22]
  wire [4:0] decode_io_decex_rsAddr_3; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_decex_rsData_0; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_decex_rsData_1; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_decex_rsData_2; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_decex_rsData_3; // @[Patmos.scala 57:22]
  wire [4:0] decode_io_decex_rdAddr_0; // @[Patmos.scala 57:22]
  wire [4:0] decode_io_decex_rdAddr_1; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_decex_immVal_0; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_decex_immVal_1; // @[Patmos.scala 57:22]
  wire  decode_io_decex_immOp_0; // @[Patmos.scala 57:22]
  wire  decode_io_decex_immOp_1; // @[Patmos.scala 57:22]
  wire  decode_io_decex_wrRd_0; // @[Patmos.scala 57:22]
  wire  decode_io_decex_wrRd_1; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_decex_callAddr; // @[Patmos.scala 57:22]
  wire  decode_io_decex_call; // @[Patmos.scala 57:22]
  wire  decode_io_decex_ret; // @[Patmos.scala 57:22]
  wire  decode_io_decex_brcf; // @[Patmos.scala 57:22]
  wire  decode_io_decex_trap; // @[Patmos.scala 57:22]
  wire  decode_io_decex_xcall; // @[Patmos.scala 57:22]
  wire  decode_io_decex_xret; // @[Patmos.scala 57:22]
  wire [4:0] decode_io_decex_xsrc; // @[Patmos.scala 57:22]
  wire  decode_io_decex_nonDelayed; // @[Patmos.scala 57:22]
  wire  decode_io_decex_illOp; // @[Patmos.scala 57:22]
  wire [4:0] decode_io_rfWrite_0_addr; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_rfWrite_0_data; // @[Patmos.scala 57:22]
  wire  decode_io_rfWrite_0_valid; // @[Patmos.scala 57:22]
  wire [4:0] decode_io_rfWrite_1_addr; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_rfWrite_1_data; // @[Patmos.scala 57:22]
  wire  decode_io_rfWrite_1_valid; // @[Patmos.scala 57:22]
  wire  decode_io_exc_exc; // @[Patmos.scala 57:22]
  wire [29:0] decode_io_exc_excBase; // @[Patmos.scala 57:22]
  wire [29:0] decode_io_exc_excAddr; // @[Patmos.scala 57:22]
  wire  decode_io_exc_intr; // @[Patmos.scala 57:22]
  wire [31:0] decode_io_exc_addr; // @[Patmos.scala 57:22]
  wire [4:0] decode_io_exc_src; // @[Patmos.scala 57:22]
  wire  decode_io_exc_local; // @[Patmos.scala 57:22]
  wire  execute_clock; // @[Patmos.scala 58:23]
  wire  execute_reset; // @[Patmos.scala 58:23]
  wire  execute_io_ena; // @[Patmos.scala 58:23]
  wire  execute_io_flush; // @[Patmos.scala 58:23]
  wire  execute_io_brflush; // @[Patmos.scala 58:23]
  wire [29:0] execute_io_decex_base; // @[Patmos.scala 58:23]
  wire [29:0] execute_io_decex_relPc; // @[Patmos.scala 58:23]
  wire [3:0] execute_io_decex_pred_0; // @[Patmos.scala 58:23]
  wire [3:0] execute_io_decex_pred_1; // @[Patmos.scala 58:23]
  wire [3:0] execute_io_decex_aluOp_0_func; // @[Patmos.scala 58:23]
  wire  execute_io_decex_aluOp_0_isMul; // @[Patmos.scala 58:23]
  wire  execute_io_decex_aluOp_0_isCmp; // @[Patmos.scala 58:23]
  wire  execute_io_decex_aluOp_0_isPred; // @[Patmos.scala 58:23]
  wire  execute_io_decex_aluOp_0_isBCpy; // @[Patmos.scala 58:23]
  wire  execute_io_decex_aluOp_0_isMTS; // @[Patmos.scala 58:23]
  wire  execute_io_decex_aluOp_0_isMFS; // @[Patmos.scala 58:23]
  wire [3:0] execute_io_decex_aluOp_1_func; // @[Patmos.scala 58:23]
  wire  execute_io_decex_aluOp_1_isCmp; // @[Patmos.scala 58:23]
  wire  execute_io_decex_aluOp_1_isPred; // @[Patmos.scala 58:23]
  wire  execute_io_decex_aluOp_1_isBCpy; // @[Patmos.scala 58:23]
  wire  execute_io_decex_aluOp_1_isMTS; // @[Patmos.scala 58:23]
  wire  execute_io_decex_aluOp_1_isMFS; // @[Patmos.scala 58:23]
  wire [1:0] execute_io_decex_predOp_0_func; // @[Patmos.scala 58:23]
  wire [2:0] execute_io_decex_predOp_0_dest; // @[Patmos.scala 58:23]
  wire [3:0] execute_io_decex_predOp_0_s1Addr; // @[Patmos.scala 58:23]
  wire [3:0] execute_io_decex_predOp_0_s2Addr; // @[Patmos.scala 58:23]
  wire [1:0] execute_io_decex_predOp_1_func; // @[Patmos.scala 58:23]
  wire [2:0] execute_io_decex_predOp_1_dest; // @[Patmos.scala 58:23]
  wire [3:0] execute_io_decex_predOp_1_s1Addr; // @[Patmos.scala 58:23]
  wire [3:0] execute_io_decex_predOp_1_s2Addr; // @[Patmos.scala 58:23]
  wire  execute_io_decex_jmpOp_branch; // @[Patmos.scala 58:23]
  wire [29:0] execute_io_decex_jmpOp_target; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_decex_jmpOp_reloc; // @[Patmos.scala 58:23]
  wire  execute_io_decex_memOp_load; // @[Patmos.scala 58:23]
  wire  execute_io_decex_memOp_store; // @[Patmos.scala 58:23]
  wire  execute_io_decex_memOp_hword; // @[Patmos.scala 58:23]
  wire  execute_io_decex_memOp_byte; // @[Patmos.scala 58:23]
  wire  execute_io_decex_memOp_zext; // @[Patmos.scala 58:23]
  wire [1:0] execute_io_decex_memOp_typ; // @[Patmos.scala 58:23]
  wire [2:0] execute_io_decex_stackOp; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_decex_rsAddr_0; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_decex_rsAddr_1; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_decex_rsAddr_2; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_decex_rsAddr_3; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_decex_rsData_0; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_decex_rsData_1; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_decex_rsData_2; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_decex_rsData_3; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_decex_rdAddr_0; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_decex_rdAddr_1; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_decex_immVal_0; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_decex_immVal_1; // @[Patmos.scala 58:23]
  wire  execute_io_decex_immOp_0; // @[Patmos.scala 58:23]
  wire  execute_io_decex_immOp_1; // @[Patmos.scala 58:23]
  wire  execute_io_decex_wrRd_0; // @[Patmos.scala 58:23]
  wire  execute_io_decex_wrRd_1; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_decex_callAddr; // @[Patmos.scala 58:23]
  wire  execute_io_decex_call; // @[Patmos.scala 58:23]
  wire  execute_io_decex_ret; // @[Patmos.scala 58:23]
  wire  execute_io_decex_brcf; // @[Patmos.scala 58:23]
  wire  execute_io_decex_trap; // @[Patmos.scala 58:23]
  wire  execute_io_decex_xcall; // @[Patmos.scala 58:23]
  wire  execute_io_decex_xret; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_decex_xsrc; // @[Patmos.scala 58:23]
  wire  execute_io_decex_nonDelayed; // @[Patmos.scala 58:23]
  wire  execute_io_decex_illOp; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_exmem_rd_0_addr; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_exmem_rd_0_data; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_rd_0_valid; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_exmem_rd_1_addr; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_exmem_rd_1_data; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_rd_1_valid; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_load; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_store; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_hword; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_byte; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_zext; // @[Patmos.scala 58:23]
  wire [1:0] execute_io_exmem_mem_typ; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_exmem_mem_addr; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_exmem_mem_data; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_call; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_ret; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_brcf; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_trap; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_xcall; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_xret; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_exmem_mem_xsrc; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_illOp; // @[Patmos.scala 58:23]
  wire  execute_io_exmem_mem_nonDelayed; // @[Patmos.scala 58:23]
  wire [29:0] execute_io_exmem_base; // @[Patmos.scala 58:23]
  wire [29:0] execute_io_exmem_relPc; // @[Patmos.scala 58:23]
  wire  execute_io_exicache_doCallRet; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_exicache_callRetBase; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_exicache_callRetAddr; // @[Patmos.scala 58:23]
  wire [29:0] execute_io_feex_pc; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_exResult_0_addr; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_exResult_0_data; // @[Patmos.scala 58:23]
  wire  execute_io_exResult_0_valid; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_exResult_1_addr; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_exResult_1_data; // @[Patmos.scala 58:23]
  wire  execute_io_exResult_1_valid; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_memResult_0_addr; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_memResult_0_data; // @[Patmos.scala 58:23]
  wire  execute_io_memResult_0_valid; // @[Patmos.scala 58:23]
  wire [4:0] execute_io_memResult_1_addr; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_memResult_1_data; // @[Patmos.scala 58:23]
  wire  execute_io_memResult_1_valid; // @[Patmos.scala 58:23]
  wire  execute_io_exfe_doBranch; // @[Patmos.scala 58:23]
  wire [29:0] execute_io_exfe_branchPc; // @[Patmos.scala 58:23]
  wire [2:0] execute_io_exsc_op; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_exsc_opData; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_exsc_opOff; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_scex_stackTop; // @[Patmos.scala 58:23]
  wire [31:0] execute_io_scex_memTop; // @[Patmos.scala 58:23]
  wire  memory_clock; // @[Patmos.scala 59:22]
  wire  memory_reset; // @[Patmos.scala 59:22]
  wire  memory_io_ena_out; // @[Patmos.scala 59:22]
  wire  memory_io_ena_in; // @[Patmos.scala 59:22]
  wire  memory_io_flush; // @[Patmos.scala 59:22]
  wire [4:0] memory_io_exmem_rd_0_addr; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_exmem_rd_0_data; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_rd_0_valid; // @[Patmos.scala 59:22]
  wire [4:0] memory_io_exmem_rd_1_addr; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_exmem_rd_1_data; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_rd_1_valid; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_load; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_store; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_hword; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_byte; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_zext; // @[Patmos.scala 59:22]
  wire [1:0] memory_io_exmem_mem_typ; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_exmem_mem_addr; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_exmem_mem_data; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_call; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_ret; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_brcf; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_trap; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_xcall; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_xret; // @[Patmos.scala 59:22]
  wire [4:0] memory_io_exmem_mem_xsrc; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_illOp; // @[Patmos.scala 59:22]
  wire  memory_io_exmem_mem_nonDelayed; // @[Patmos.scala 59:22]
  wire [29:0] memory_io_exmem_base; // @[Patmos.scala 59:22]
  wire [29:0] memory_io_exmem_relPc; // @[Patmos.scala 59:22]
  wire [4:0] memory_io_memwb_rd_0_addr; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_memwb_rd_0_data; // @[Patmos.scala 59:22]
  wire  memory_io_memwb_rd_0_valid; // @[Patmos.scala 59:22]
  wire [4:0] memory_io_memwb_rd_1_addr; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_memwb_rd_1_data; // @[Patmos.scala 59:22]
  wire  memory_io_memwb_rd_1_valid; // @[Patmos.scala 59:22]
  wire  memory_io_memfe_doCallRet; // @[Patmos.scala 59:22]
  wire  memory_io_memfe_store; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_memfe_addr; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_memfe_data; // @[Patmos.scala 59:22]
  wire [4:0] memory_io_exResult_0_addr; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_exResult_0_data; // @[Patmos.scala 59:22]
  wire  memory_io_exResult_0_valid; // @[Patmos.scala 59:22]
  wire [4:0] memory_io_exResult_1_addr; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_exResult_1_data; // @[Patmos.scala 59:22]
  wire  memory_io_exResult_1_valid; // @[Patmos.scala 59:22]
  wire [2:0] memory_io_localInOut_M_Cmd; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_localInOut_M_Addr; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_localInOut_M_Data; // @[Patmos.scala 59:22]
  wire [3:0] memory_io_localInOut_M_ByteEn; // @[Patmos.scala 59:22]
  wire [1:0] memory_io_localInOut_S_Resp; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_localInOut_S_Data; // @[Patmos.scala 59:22]
  wire [2:0] memory_io_globalInOut_M_Cmd; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_globalInOut_M_Addr; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_globalInOut_M_Data; // @[Patmos.scala 59:22]
  wire [3:0] memory_io_globalInOut_M_ByteEn; // @[Patmos.scala 59:22]
  wire [1:0] memory_io_globalInOut_M_AddrSpace; // @[Patmos.scala 59:22]
  wire [1:0] memory_io_globalInOut_S_Resp; // @[Patmos.scala 59:22]
  wire [31:0] memory_io_globalInOut_S_Data; // @[Patmos.scala 59:22]
  wire  memory_io_icacheIllMem; // @[Patmos.scala 59:22]
  wire  memory_io_scacheIllMem; // @[Patmos.scala 59:22]
  wire  memory_io_exc_call; // @[Patmos.scala 59:22]
  wire  memory_io_exc_ret; // @[Patmos.scala 59:22]
  wire [4:0] memory_io_exc_src; // @[Patmos.scala 59:22]
  wire  memory_io_exc_exc; // @[Patmos.scala 59:22]
  wire [29:0] memory_io_exc_excBase; // @[Patmos.scala 59:22]
  wire [29:0] memory_io_exc_excAddr; // @[Patmos.scala 59:22]
  wire [4:0] writeback_io_memwb_rd_0_addr; // @[Patmos.scala 60:25]
  wire [31:0] writeback_io_memwb_rd_0_data; // @[Patmos.scala 60:25]
  wire  writeback_io_memwb_rd_0_valid; // @[Patmos.scala 60:25]
  wire [4:0] writeback_io_memwb_rd_1_addr; // @[Patmos.scala 60:25]
  wire [31:0] writeback_io_memwb_rd_1_data; // @[Patmos.scala 60:25]
  wire  writeback_io_memwb_rd_1_valid; // @[Patmos.scala 60:25]
  wire [4:0] writeback_io_rfWrite_0_addr; // @[Patmos.scala 60:25]
  wire [31:0] writeback_io_rfWrite_0_data; // @[Patmos.scala 60:25]
  wire  writeback_io_rfWrite_0_valid; // @[Patmos.scala 60:25]
  wire [4:0] writeback_io_rfWrite_1_addr; // @[Patmos.scala 60:25]
  wire [31:0] writeback_io_rfWrite_1_data; // @[Patmos.scala 60:25]
  wire  writeback_io_rfWrite_1_valid; // @[Patmos.scala 60:25]
  wire [4:0] writeback_io_memResult_0_addr; // @[Patmos.scala 60:25]
  wire [31:0] writeback_io_memResult_0_data; // @[Patmos.scala 60:25]
  wire  writeback_io_memResult_0_valid; // @[Patmos.scala 60:25]
  wire [4:0] writeback_io_memResult_1_addr; // @[Patmos.scala 60:25]
  wire [31:0] writeback_io_memResult_1_data; // @[Patmos.scala 60:25]
  wire  writeback_io_memResult_1_valid; // @[Patmos.scala 60:25]
  wire  exc_clock; // @[Patmos.scala 61:19]
  wire  exc_reset; // @[Patmos.scala 61:19]
  wire  exc_io_ena; // @[Patmos.scala 61:19]
  wire [2:0] exc_io_ocp_M_Cmd; // @[Patmos.scala 61:19]
  wire [31:0] exc_io_ocp_M_Addr; // @[Patmos.scala 61:19]
  wire [31:0] exc_io_ocp_M_Data; // @[Patmos.scala 61:19]
  wire [1:0] exc_io_ocp_S_Resp; // @[Patmos.scala 61:19]
  wire [31:0] exc_io_ocp_S_Data; // @[Patmos.scala 61:19]
  wire  exc_io_intrs_0; // @[Patmos.scala 61:19]
  wire  exc_io_intrs_1; // @[Patmos.scala 61:19]
  wire  exc_io_intrs_2; // @[Patmos.scala 61:19]
  wire  exc_io_intrs_3; // @[Patmos.scala 61:19]
  wire  exc_io_intrs_4; // @[Patmos.scala 61:19]
  wire  exc_io_intrs_5; // @[Patmos.scala 61:19]
  wire  exc_io_excdec_exc; // @[Patmos.scala 61:19]
  wire [29:0] exc_io_excdec_excBase; // @[Patmos.scala 61:19]
  wire [29:0] exc_io_excdec_excAddr; // @[Patmos.scala 61:19]
  wire  exc_io_excdec_intr; // @[Patmos.scala 61:19]
  wire [31:0] exc_io_excdec_addr; // @[Patmos.scala 61:19]
  wire [4:0] exc_io_excdec_src; // @[Patmos.scala 61:19]
  wire  exc_io_excdec_local; // @[Patmos.scala 61:19]
  wire  exc_io_memexc_call; // @[Patmos.scala 61:19]
  wire  exc_io_memexc_ret; // @[Patmos.scala 61:19]
  wire [4:0] exc_io_memexc_src; // @[Patmos.scala 61:19]
  wire  exc_io_memexc_exc; // @[Patmos.scala 61:19]
  wire [29:0] exc_io_memexc_excBase; // @[Patmos.scala 61:19]
  wire [29:0] exc_io_memexc_excAddr; // @[Patmos.scala 61:19]
  wire  exc_io_invalICache; // @[Patmos.scala 61:19]
  wire  exc_io_invalDCache; // @[Patmos.scala 61:19]
  wire  dcache_clock; // @[Patmos.scala 63:22]
  wire  dcache_reset; // @[Patmos.scala 63:22]
  wire [2:0] dcache_io_master_M_Cmd; // @[Patmos.scala 63:22]
  wire [31:0] dcache_io_master_M_Addr; // @[Patmos.scala 63:22]
  wire [31:0] dcache_io_master_M_Data; // @[Patmos.scala 63:22]
  wire [3:0] dcache_io_master_M_ByteEn; // @[Patmos.scala 63:22]
  wire [1:0] dcache_io_master_M_AddrSpace; // @[Patmos.scala 63:22]
  wire [1:0] dcache_io_master_S_Resp; // @[Patmos.scala 63:22]
  wire [31:0] dcache_io_master_S_Data; // @[Patmos.scala 63:22]
  wire [2:0] dcache_io_slave_M_Cmd; // @[Patmos.scala 63:22]
  wire [31:0] dcache_io_slave_M_Addr; // @[Patmos.scala 63:22]
  wire [31:0] dcache_io_slave_M_Data; // @[Patmos.scala 63:22]
  wire  dcache_io_slave_M_DataValid; // @[Patmos.scala 63:22]
  wire [3:0] dcache_io_slave_M_DataByteEn; // @[Patmos.scala 63:22]
  wire [1:0] dcache_io_slave_S_Resp; // @[Patmos.scala 63:22]
  wire [31:0] dcache_io_slave_S_Data; // @[Patmos.scala 63:22]
  wire  dcache_io_slave_S_CmdAccept; // @[Patmos.scala 63:22]
  wire  dcache_io_slave_S_DataAccept; // @[Patmos.scala 63:22]
  wire  dcache_io_scIO_ena_in; // @[Patmos.scala 63:22]
  wire [2:0] dcache_io_scIO_exsc_op; // @[Patmos.scala 63:22]
  wire [31:0] dcache_io_scIO_exsc_opData; // @[Patmos.scala 63:22]
  wire [31:0] dcache_io_scIO_exsc_opOff; // @[Patmos.scala 63:22]
  wire [31:0] dcache_io_scIO_scex_stackTop; // @[Patmos.scala 63:22]
  wire [31:0] dcache_io_scIO_scex_memTop; // @[Patmos.scala 63:22]
  wire  dcache_io_scIO_illMem; // @[Patmos.scala 63:22]
  wire  dcache_io_scIO_stall; // @[Patmos.scala 63:22]
  wire  dcache_io_invalDCache; // @[Patmos.scala 63:22]
  wire [2:0] burstBus_io_master_M_Cmd; // @[Patmos.scala 107:24]
  wire [31:0] burstBus_io_master_M_Addr; // @[Patmos.scala 107:24]
  wire [31:0] burstBus_io_master_M_Data; // @[Patmos.scala 107:24]
  wire  burstBus_io_master_M_DataValid; // @[Patmos.scala 107:24]
  wire [3:0] burstBus_io_master_M_DataByteEn; // @[Patmos.scala 107:24]
  wire [1:0] burstBus_io_master_S_Resp; // @[Patmos.scala 107:24]
  wire [31:0] burstBus_io_master_S_Data; // @[Patmos.scala 107:24]
  wire  burstBus_io_master_S_CmdAccept; // @[Patmos.scala 107:24]
  wire  burstBus_io_master_S_DataAccept; // @[Patmos.scala 107:24]
  wire [2:0] burstBus_io_slave_M_Cmd; // @[Patmos.scala 107:24]
  wire [31:0] burstBus_io_slave_M_Addr; // @[Patmos.scala 107:24]
  wire [31:0] burstBus_io_slave_M_Data; // @[Patmos.scala 107:24]
  wire  burstBus_io_slave_M_DataValid; // @[Patmos.scala 107:24]
  wire [3:0] burstBus_io_slave_M_DataByteEn; // @[Patmos.scala 107:24]
  wire [1:0] burstBus_io_slave_S_Resp; // @[Patmos.scala 107:24]
  wire [31:0] burstBus_io_slave_S_Data; // @[Patmos.scala 107:24]
  wire  burstBus_io_slave_S_CmdAccept; // @[Patmos.scala 107:24]
  wire  burstBus_io_slave_S_DataAccept; // @[Patmos.scala 107:24]
  wire [2:0] mmu_io_virt_M_Cmd; // @[Patmos.scala 119:19]
  wire [31:0] mmu_io_virt_M_Addr; // @[Patmos.scala 119:19]
  wire [31:0] mmu_io_virt_M_Data; // @[Patmos.scala 119:19]
  wire  mmu_io_virt_M_DataValid; // @[Patmos.scala 119:19]
  wire [3:0] mmu_io_virt_M_DataByteEn; // @[Patmos.scala 119:19]
  wire [1:0] mmu_io_virt_S_Resp; // @[Patmos.scala 119:19]
  wire [31:0] mmu_io_virt_S_Data; // @[Patmos.scala 119:19]
  wire [2:0] mmu_io_phys_M_Cmd; // @[Patmos.scala 119:19]
  wire [20:0] mmu_io_phys_M_Addr; // @[Patmos.scala 119:19]
  wire [31:0] mmu_io_phys_M_Data; // @[Patmos.scala 119:19]
  wire  mmu_io_phys_M_DataValid; // @[Patmos.scala 119:19]
  wire [3:0] mmu_io_phys_M_DataByteEn; // @[Patmos.scala 119:19]
  wire [1:0] mmu_io_phys_S_Resp; // @[Patmos.scala 119:19]
  wire [31:0] mmu_io_phys_S_Data; // @[Patmos.scala 119:19]
  reg  REG; // @[OcpBurst.scala 144:24]
  wire  _T_2 = dcache_io_slave_M_Cmd != 3'h0 | REG; // @[OcpBurst.scala 147:25]
  wire  _T_3 = icache_io_ocp_port_M_Cmd != 3'h0 ? 1'h0 : _T_2; // @[OcpBurst.scala 146:18]
  wire  _T_6 = ~dcache_io_scIO_stall; // @[Patmos.scala 126:44]
  wire  _T_10 = memory_io_ena_out & icache_io_ena_out; // @[Patmos.scala 128:46]
  reg  enableReg; // @[Patmos.scala 137:22]
  MCache icache ( // @[Patmos.scala 44:13]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_ena_out(icache_io_ena_out),
    .io_ena_in(icache_io_ena_in),
    .io_invalidate(icache_io_invalidate),
    .io_feicache_addrEven(icache_io_feicache_addrEven),
    .io_feicache_addrOdd(icache_io_feicache_addrOdd),
    .io_exicache_doCallRet(icache_io_exicache_doCallRet),
    .io_exicache_callRetBase(icache_io_exicache_callRetBase),
    .io_exicache_callRetAddr(icache_io_exicache_callRetAddr),
    .io_icachefe_instrEven(icache_io_icachefe_instrEven),
    .io_icachefe_instrOdd(icache_io_icachefe_instrOdd),
    .io_icachefe_base(icache_io_icachefe_base),
    .io_icachefe_relBase(icache_io_icachefe_relBase),
    .io_icachefe_relPc(icache_io_icachefe_relPc),
    .io_icachefe_reloc(icache_io_icachefe_reloc),
    .io_icachefe_memSel(icache_io_icachefe_memSel),
    .io_ocp_port_M_Cmd(icache_io_ocp_port_M_Cmd),
    .io_ocp_port_M_Addr(icache_io_ocp_port_M_Addr),
    .io_ocp_port_S_Resp(icache_io_ocp_port_S_Resp),
    .io_ocp_port_S_Data(icache_io_ocp_port_S_Data),
    .io_ocp_port_S_CmdAccept(icache_io_ocp_port_S_CmdAccept),
    .io_illMem(icache_io_illMem)
  );
  Fetch fetch ( // @[Patmos.scala 56:21]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_ena(fetch_io_ena),
    .io_fedec_instr_a(fetch_io_fedec_instr_a),
    .io_fedec_instr_b(fetch_io_fedec_instr_b),
    .io_fedec_pc(fetch_io_fedec_pc),
    .io_fedec_base(fetch_io_fedec_base),
    .io_fedec_reloc(fetch_io_fedec_reloc),
    .io_fedec_relPc(fetch_io_fedec_relPc),
    .io_feex_pc(fetch_io_feex_pc),
    .io_exfe_doBranch(fetch_io_exfe_doBranch),
    .io_exfe_branchPc(fetch_io_exfe_branchPc),
    .io_memfe_doCallRet(fetch_io_memfe_doCallRet),
    .io_memfe_store(fetch_io_memfe_store),
    .io_memfe_addr(fetch_io_memfe_addr),
    .io_memfe_data(fetch_io_memfe_data),
    .io_feicache_addrEven(fetch_io_feicache_addrEven),
    .io_feicache_addrOdd(fetch_io_feicache_addrOdd),
    .io_icachefe_instrEven(fetch_io_icachefe_instrEven),
    .io_icachefe_instrOdd(fetch_io_icachefe_instrOdd),
    .io_icachefe_base(fetch_io_icachefe_base),
    .io_icachefe_relBase(fetch_io_icachefe_relBase),
    .io_icachefe_relPc(fetch_io_icachefe_relPc),
    .io_icachefe_reloc(fetch_io_icachefe_reloc),
    .io_icachefe_memSel(fetch_io_icachefe_memSel)
  );
  Decode decode ( // @[Patmos.scala 57:22]
    .clock(decode_clock),
    .reset(decode_reset),
    .io_ena(decode_io_ena),
    .io_flush(decode_io_flush),
    .io_fedec_instr_a(decode_io_fedec_instr_a),
    .io_fedec_instr_b(decode_io_fedec_instr_b),
    .io_fedec_pc(decode_io_fedec_pc),
    .io_fedec_base(decode_io_fedec_base),
    .io_fedec_reloc(decode_io_fedec_reloc),
    .io_fedec_relPc(decode_io_fedec_relPc),
    .io_decex_base(decode_io_decex_base),
    .io_decex_relPc(decode_io_decex_relPc),
    .io_decex_pred_0(decode_io_decex_pred_0),
    .io_decex_pred_1(decode_io_decex_pred_1),
    .io_decex_aluOp_0_func(decode_io_decex_aluOp_0_func),
    .io_decex_aluOp_0_isMul(decode_io_decex_aluOp_0_isMul),
    .io_decex_aluOp_0_isCmp(decode_io_decex_aluOp_0_isCmp),
    .io_decex_aluOp_0_isPred(decode_io_decex_aluOp_0_isPred),
    .io_decex_aluOp_0_isBCpy(decode_io_decex_aluOp_0_isBCpy),
    .io_decex_aluOp_0_isMTS(decode_io_decex_aluOp_0_isMTS),
    .io_decex_aluOp_0_isMFS(decode_io_decex_aluOp_0_isMFS),
    .io_decex_aluOp_1_func(decode_io_decex_aluOp_1_func),
    .io_decex_aluOp_1_isCmp(decode_io_decex_aluOp_1_isCmp),
    .io_decex_aluOp_1_isPred(decode_io_decex_aluOp_1_isPred),
    .io_decex_aluOp_1_isBCpy(decode_io_decex_aluOp_1_isBCpy),
    .io_decex_aluOp_1_isMTS(decode_io_decex_aluOp_1_isMTS),
    .io_decex_aluOp_1_isMFS(decode_io_decex_aluOp_1_isMFS),
    .io_decex_predOp_0_func(decode_io_decex_predOp_0_func),
    .io_decex_predOp_0_dest(decode_io_decex_predOp_0_dest),
    .io_decex_predOp_0_s1Addr(decode_io_decex_predOp_0_s1Addr),
    .io_decex_predOp_0_s2Addr(decode_io_decex_predOp_0_s2Addr),
    .io_decex_predOp_1_func(decode_io_decex_predOp_1_func),
    .io_decex_predOp_1_dest(decode_io_decex_predOp_1_dest),
    .io_decex_predOp_1_s1Addr(decode_io_decex_predOp_1_s1Addr),
    .io_decex_predOp_1_s2Addr(decode_io_decex_predOp_1_s2Addr),
    .io_decex_jmpOp_branch(decode_io_decex_jmpOp_branch),
    .io_decex_jmpOp_target(decode_io_decex_jmpOp_target),
    .io_decex_jmpOp_reloc(decode_io_decex_jmpOp_reloc),
    .io_decex_memOp_load(decode_io_decex_memOp_load),
    .io_decex_memOp_store(decode_io_decex_memOp_store),
    .io_decex_memOp_hword(decode_io_decex_memOp_hword),
    .io_decex_memOp_byte(decode_io_decex_memOp_byte),
    .io_decex_memOp_zext(decode_io_decex_memOp_zext),
    .io_decex_memOp_typ(decode_io_decex_memOp_typ),
    .io_decex_stackOp(decode_io_decex_stackOp),
    .io_decex_rsAddr_0(decode_io_decex_rsAddr_0),
    .io_decex_rsAddr_1(decode_io_decex_rsAddr_1),
    .io_decex_rsAddr_2(decode_io_decex_rsAddr_2),
    .io_decex_rsAddr_3(decode_io_decex_rsAddr_3),
    .io_decex_rsData_0(decode_io_decex_rsData_0),
    .io_decex_rsData_1(decode_io_decex_rsData_1),
    .io_decex_rsData_2(decode_io_decex_rsData_2),
    .io_decex_rsData_3(decode_io_decex_rsData_3),
    .io_decex_rdAddr_0(decode_io_decex_rdAddr_0),
    .io_decex_rdAddr_1(decode_io_decex_rdAddr_1),
    .io_decex_immVal_0(decode_io_decex_immVal_0),
    .io_decex_immVal_1(decode_io_decex_immVal_1),
    .io_decex_immOp_0(decode_io_decex_immOp_0),
    .io_decex_immOp_1(decode_io_decex_immOp_1),
    .io_decex_wrRd_0(decode_io_decex_wrRd_0),
    .io_decex_wrRd_1(decode_io_decex_wrRd_1),
    .io_decex_callAddr(decode_io_decex_callAddr),
    .io_decex_call(decode_io_decex_call),
    .io_decex_ret(decode_io_decex_ret),
    .io_decex_brcf(decode_io_decex_brcf),
    .io_decex_trap(decode_io_decex_trap),
    .io_decex_xcall(decode_io_decex_xcall),
    .io_decex_xret(decode_io_decex_xret),
    .io_decex_xsrc(decode_io_decex_xsrc),
    .io_decex_nonDelayed(decode_io_decex_nonDelayed),
    .io_decex_illOp(decode_io_decex_illOp),
    .io_rfWrite_0_addr(decode_io_rfWrite_0_addr),
    .io_rfWrite_0_data(decode_io_rfWrite_0_data),
    .io_rfWrite_0_valid(decode_io_rfWrite_0_valid),
    .io_rfWrite_1_addr(decode_io_rfWrite_1_addr),
    .io_rfWrite_1_data(decode_io_rfWrite_1_data),
    .io_rfWrite_1_valid(decode_io_rfWrite_1_valid),
    .io_exc_exc(decode_io_exc_exc),
    .io_exc_excBase(decode_io_exc_excBase),
    .io_exc_excAddr(decode_io_exc_excAddr),
    .io_exc_intr(decode_io_exc_intr),
    .io_exc_addr(decode_io_exc_addr),
    .io_exc_src(decode_io_exc_src),
    .io_exc_local(decode_io_exc_local)
  );
  Execute execute ( // @[Patmos.scala 58:23]
    .clock(execute_clock),
    .reset(execute_reset),
    .io_ena(execute_io_ena),
    .io_flush(execute_io_flush),
    .io_brflush(execute_io_brflush),
    .io_decex_base(execute_io_decex_base),
    .io_decex_relPc(execute_io_decex_relPc),
    .io_decex_pred_0(execute_io_decex_pred_0),
    .io_decex_pred_1(execute_io_decex_pred_1),
    .io_decex_aluOp_0_func(execute_io_decex_aluOp_0_func),
    .io_decex_aluOp_0_isMul(execute_io_decex_aluOp_0_isMul),
    .io_decex_aluOp_0_isCmp(execute_io_decex_aluOp_0_isCmp),
    .io_decex_aluOp_0_isPred(execute_io_decex_aluOp_0_isPred),
    .io_decex_aluOp_0_isBCpy(execute_io_decex_aluOp_0_isBCpy),
    .io_decex_aluOp_0_isMTS(execute_io_decex_aluOp_0_isMTS),
    .io_decex_aluOp_0_isMFS(execute_io_decex_aluOp_0_isMFS),
    .io_decex_aluOp_1_func(execute_io_decex_aluOp_1_func),
    .io_decex_aluOp_1_isCmp(execute_io_decex_aluOp_1_isCmp),
    .io_decex_aluOp_1_isPred(execute_io_decex_aluOp_1_isPred),
    .io_decex_aluOp_1_isBCpy(execute_io_decex_aluOp_1_isBCpy),
    .io_decex_aluOp_1_isMTS(execute_io_decex_aluOp_1_isMTS),
    .io_decex_aluOp_1_isMFS(execute_io_decex_aluOp_1_isMFS),
    .io_decex_predOp_0_func(execute_io_decex_predOp_0_func),
    .io_decex_predOp_0_dest(execute_io_decex_predOp_0_dest),
    .io_decex_predOp_0_s1Addr(execute_io_decex_predOp_0_s1Addr),
    .io_decex_predOp_0_s2Addr(execute_io_decex_predOp_0_s2Addr),
    .io_decex_predOp_1_func(execute_io_decex_predOp_1_func),
    .io_decex_predOp_1_dest(execute_io_decex_predOp_1_dest),
    .io_decex_predOp_1_s1Addr(execute_io_decex_predOp_1_s1Addr),
    .io_decex_predOp_1_s2Addr(execute_io_decex_predOp_1_s2Addr),
    .io_decex_jmpOp_branch(execute_io_decex_jmpOp_branch),
    .io_decex_jmpOp_target(execute_io_decex_jmpOp_target),
    .io_decex_jmpOp_reloc(execute_io_decex_jmpOp_reloc),
    .io_decex_memOp_load(execute_io_decex_memOp_load),
    .io_decex_memOp_store(execute_io_decex_memOp_store),
    .io_decex_memOp_hword(execute_io_decex_memOp_hword),
    .io_decex_memOp_byte(execute_io_decex_memOp_byte),
    .io_decex_memOp_zext(execute_io_decex_memOp_zext),
    .io_decex_memOp_typ(execute_io_decex_memOp_typ),
    .io_decex_stackOp(execute_io_decex_stackOp),
    .io_decex_rsAddr_0(execute_io_decex_rsAddr_0),
    .io_decex_rsAddr_1(execute_io_decex_rsAddr_1),
    .io_decex_rsAddr_2(execute_io_decex_rsAddr_2),
    .io_decex_rsAddr_3(execute_io_decex_rsAddr_3),
    .io_decex_rsData_0(execute_io_decex_rsData_0),
    .io_decex_rsData_1(execute_io_decex_rsData_1),
    .io_decex_rsData_2(execute_io_decex_rsData_2),
    .io_decex_rsData_3(execute_io_decex_rsData_3),
    .io_decex_rdAddr_0(execute_io_decex_rdAddr_0),
    .io_decex_rdAddr_1(execute_io_decex_rdAddr_1),
    .io_decex_immVal_0(execute_io_decex_immVal_0),
    .io_decex_immVal_1(execute_io_decex_immVal_1),
    .io_decex_immOp_0(execute_io_decex_immOp_0),
    .io_decex_immOp_1(execute_io_decex_immOp_1),
    .io_decex_wrRd_0(execute_io_decex_wrRd_0),
    .io_decex_wrRd_1(execute_io_decex_wrRd_1),
    .io_decex_callAddr(execute_io_decex_callAddr),
    .io_decex_call(execute_io_decex_call),
    .io_decex_ret(execute_io_decex_ret),
    .io_decex_brcf(execute_io_decex_brcf),
    .io_decex_trap(execute_io_decex_trap),
    .io_decex_xcall(execute_io_decex_xcall),
    .io_decex_xret(execute_io_decex_xret),
    .io_decex_xsrc(execute_io_decex_xsrc),
    .io_decex_nonDelayed(execute_io_decex_nonDelayed),
    .io_decex_illOp(execute_io_decex_illOp),
    .io_exmem_rd_0_addr(execute_io_exmem_rd_0_addr),
    .io_exmem_rd_0_data(execute_io_exmem_rd_0_data),
    .io_exmem_rd_0_valid(execute_io_exmem_rd_0_valid),
    .io_exmem_rd_1_addr(execute_io_exmem_rd_1_addr),
    .io_exmem_rd_1_data(execute_io_exmem_rd_1_data),
    .io_exmem_rd_1_valid(execute_io_exmem_rd_1_valid),
    .io_exmem_mem_load(execute_io_exmem_mem_load),
    .io_exmem_mem_store(execute_io_exmem_mem_store),
    .io_exmem_mem_hword(execute_io_exmem_mem_hword),
    .io_exmem_mem_byte(execute_io_exmem_mem_byte),
    .io_exmem_mem_zext(execute_io_exmem_mem_zext),
    .io_exmem_mem_typ(execute_io_exmem_mem_typ),
    .io_exmem_mem_addr(execute_io_exmem_mem_addr),
    .io_exmem_mem_data(execute_io_exmem_mem_data),
    .io_exmem_mem_call(execute_io_exmem_mem_call),
    .io_exmem_mem_ret(execute_io_exmem_mem_ret),
    .io_exmem_mem_brcf(execute_io_exmem_mem_brcf),
    .io_exmem_mem_trap(execute_io_exmem_mem_trap),
    .io_exmem_mem_xcall(execute_io_exmem_mem_xcall),
    .io_exmem_mem_xret(execute_io_exmem_mem_xret),
    .io_exmem_mem_xsrc(execute_io_exmem_mem_xsrc),
    .io_exmem_mem_illOp(execute_io_exmem_mem_illOp),
    .io_exmem_mem_nonDelayed(execute_io_exmem_mem_nonDelayed),
    .io_exmem_base(execute_io_exmem_base),
    .io_exmem_relPc(execute_io_exmem_relPc),
    .io_exicache_doCallRet(execute_io_exicache_doCallRet),
    .io_exicache_callRetBase(execute_io_exicache_callRetBase),
    .io_exicache_callRetAddr(execute_io_exicache_callRetAddr),
    .io_feex_pc(execute_io_feex_pc),
    .io_exResult_0_addr(execute_io_exResult_0_addr),
    .io_exResult_0_data(execute_io_exResult_0_data),
    .io_exResult_0_valid(execute_io_exResult_0_valid),
    .io_exResult_1_addr(execute_io_exResult_1_addr),
    .io_exResult_1_data(execute_io_exResult_1_data),
    .io_exResult_1_valid(execute_io_exResult_1_valid),
    .io_memResult_0_addr(execute_io_memResult_0_addr),
    .io_memResult_0_data(execute_io_memResult_0_data),
    .io_memResult_0_valid(execute_io_memResult_0_valid),
    .io_memResult_1_addr(execute_io_memResult_1_addr),
    .io_memResult_1_data(execute_io_memResult_1_data),
    .io_memResult_1_valid(execute_io_memResult_1_valid),
    .io_exfe_doBranch(execute_io_exfe_doBranch),
    .io_exfe_branchPc(execute_io_exfe_branchPc),
    .io_exsc_op(execute_io_exsc_op),
    .io_exsc_opData(execute_io_exsc_opData),
    .io_exsc_opOff(execute_io_exsc_opOff),
    .io_scex_stackTop(execute_io_scex_stackTop),
    .io_scex_memTop(execute_io_scex_memTop)
  );
  Memory memory ( // @[Patmos.scala 59:22]
    .clock(memory_clock),
    .reset(memory_reset),
    .io_ena_out(memory_io_ena_out),
    .io_ena_in(memory_io_ena_in),
    .io_flush(memory_io_flush),
    .io_exmem_rd_0_addr(memory_io_exmem_rd_0_addr),
    .io_exmem_rd_0_data(memory_io_exmem_rd_0_data),
    .io_exmem_rd_0_valid(memory_io_exmem_rd_0_valid),
    .io_exmem_rd_1_addr(memory_io_exmem_rd_1_addr),
    .io_exmem_rd_1_data(memory_io_exmem_rd_1_data),
    .io_exmem_rd_1_valid(memory_io_exmem_rd_1_valid),
    .io_exmem_mem_load(memory_io_exmem_mem_load),
    .io_exmem_mem_store(memory_io_exmem_mem_store),
    .io_exmem_mem_hword(memory_io_exmem_mem_hword),
    .io_exmem_mem_byte(memory_io_exmem_mem_byte),
    .io_exmem_mem_zext(memory_io_exmem_mem_zext),
    .io_exmem_mem_typ(memory_io_exmem_mem_typ),
    .io_exmem_mem_addr(memory_io_exmem_mem_addr),
    .io_exmem_mem_data(memory_io_exmem_mem_data),
    .io_exmem_mem_call(memory_io_exmem_mem_call),
    .io_exmem_mem_ret(memory_io_exmem_mem_ret),
    .io_exmem_mem_brcf(memory_io_exmem_mem_brcf),
    .io_exmem_mem_trap(memory_io_exmem_mem_trap),
    .io_exmem_mem_xcall(memory_io_exmem_mem_xcall),
    .io_exmem_mem_xret(memory_io_exmem_mem_xret),
    .io_exmem_mem_xsrc(memory_io_exmem_mem_xsrc),
    .io_exmem_mem_illOp(memory_io_exmem_mem_illOp),
    .io_exmem_mem_nonDelayed(memory_io_exmem_mem_nonDelayed),
    .io_exmem_base(memory_io_exmem_base),
    .io_exmem_relPc(memory_io_exmem_relPc),
    .io_memwb_rd_0_addr(memory_io_memwb_rd_0_addr),
    .io_memwb_rd_0_data(memory_io_memwb_rd_0_data),
    .io_memwb_rd_0_valid(memory_io_memwb_rd_0_valid),
    .io_memwb_rd_1_addr(memory_io_memwb_rd_1_addr),
    .io_memwb_rd_1_data(memory_io_memwb_rd_1_data),
    .io_memwb_rd_1_valid(memory_io_memwb_rd_1_valid),
    .io_memfe_doCallRet(memory_io_memfe_doCallRet),
    .io_memfe_store(memory_io_memfe_store),
    .io_memfe_addr(memory_io_memfe_addr),
    .io_memfe_data(memory_io_memfe_data),
    .io_exResult_0_addr(memory_io_exResult_0_addr),
    .io_exResult_0_data(memory_io_exResult_0_data),
    .io_exResult_0_valid(memory_io_exResult_0_valid),
    .io_exResult_1_addr(memory_io_exResult_1_addr),
    .io_exResult_1_data(memory_io_exResult_1_data),
    .io_exResult_1_valid(memory_io_exResult_1_valid),
    .io_localInOut_M_Cmd(memory_io_localInOut_M_Cmd),
    .io_localInOut_M_Addr(memory_io_localInOut_M_Addr),
    .io_localInOut_M_Data(memory_io_localInOut_M_Data),
    .io_localInOut_M_ByteEn(memory_io_localInOut_M_ByteEn),
    .io_localInOut_S_Resp(memory_io_localInOut_S_Resp),
    .io_localInOut_S_Data(memory_io_localInOut_S_Data),
    .io_globalInOut_M_Cmd(memory_io_globalInOut_M_Cmd),
    .io_globalInOut_M_Addr(memory_io_globalInOut_M_Addr),
    .io_globalInOut_M_Data(memory_io_globalInOut_M_Data),
    .io_globalInOut_M_ByteEn(memory_io_globalInOut_M_ByteEn),
    .io_globalInOut_M_AddrSpace(memory_io_globalInOut_M_AddrSpace),
    .io_globalInOut_S_Resp(memory_io_globalInOut_S_Resp),
    .io_globalInOut_S_Data(memory_io_globalInOut_S_Data),
    .io_icacheIllMem(memory_io_icacheIllMem),
    .io_scacheIllMem(memory_io_scacheIllMem),
    .io_exc_call(memory_io_exc_call),
    .io_exc_ret(memory_io_exc_ret),
    .io_exc_src(memory_io_exc_src),
    .io_exc_exc(memory_io_exc_exc),
    .io_exc_excBase(memory_io_exc_excBase),
    .io_exc_excAddr(memory_io_exc_excAddr)
  );
  WriteBack writeback ( // @[Patmos.scala 60:25]
    .io_memwb_rd_0_addr(writeback_io_memwb_rd_0_addr),
    .io_memwb_rd_0_data(writeback_io_memwb_rd_0_data),
    .io_memwb_rd_0_valid(writeback_io_memwb_rd_0_valid),
    .io_memwb_rd_1_addr(writeback_io_memwb_rd_1_addr),
    .io_memwb_rd_1_data(writeback_io_memwb_rd_1_data),
    .io_memwb_rd_1_valid(writeback_io_memwb_rd_1_valid),
    .io_rfWrite_0_addr(writeback_io_rfWrite_0_addr),
    .io_rfWrite_0_data(writeback_io_rfWrite_0_data),
    .io_rfWrite_0_valid(writeback_io_rfWrite_0_valid),
    .io_rfWrite_1_addr(writeback_io_rfWrite_1_addr),
    .io_rfWrite_1_data(writeback_io_rfWrite_1_data),
    .io_rfWrite_1_valid(writeback_io_rfWrite_1_valid),
    .io_memResult_0_addr(writeback_io_memResult_0_addr),
    .io_memResult_0_data(writeback_io_memResult_0_data),
    .io_memResult_0_valid(writeback_io_memResult_0_valid),
    .io_memResult_1_addr(writeback_io_memResult_1_addr),
    .io_memResult_1_data(writeback_io_memResult_1_data),
    .io_memResult_1_valid(writeback_io_memResult_1_valid)
  );
  Exceptions exc ( // @[Patmos.scala 61:19]
    .clock(exc_clock),
    .reset(exc_reset),
    .io_ena(exc_io_ena),
    .io_ocp_M_Cmd(exc_io_ocp_M_Cmd),
    .io_ocp_M_Addr(exc_io_ocp_M_Addr),
    .io_ocp_M_Data(exc_io_ocp_M_Data),
    .io_ocp_S_Resp(exc_io_ocp_S_Resp),
    .io_ocp_S_Data(exc_io_ocp_S_Data),
    .io_intrs_0(exc_io_intrs_0),
    .io_intrs_1(exc_io_intrs_1),
    .io_intrs_2(exc_io_intrs_2),
    .io_intrs_3(exc_io_intrs_3),
    .io_intrs_4(exc_io_intrs_4),
    .io_intrs_5(exc_io_intrs_5),
    .io_excdec_exc(exc_io_excdec_exc),
    .io_excdec_excBase(exc_io_excdec_excBase),
    .io_excdec_excAddr(exc_io_excdec_excAddr),
    .io_excdec_intr(exc_io_excdec_intr),
    .io_excdec_addr(exc_io_excdec_addr),
    .io_excdec_src(exc_io_excdec_src),
    .io_excdec_local(exc_io_excdec_local),
    .io_memexc_call(exc_io_memexc_call),
    .io_memexc_ret(exc_io_memexc_ret),
    .io_memexc_src(exc_io_memexc_src),
    .io_memexc_exc(exc_io_memexc_exc),
    .io_memexc_excBase(exc_io_memexc_excBase),
    .io_memexc_excAddr(exc_io_memexc_excAddr),
    .io_invalICache(exc_io_invalICache),
    .io_invalDCache(exc_io_invalDCache)
  );
  DataCache dcache ( // @[Patmos.scala 63:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_master_M_Cmd(dcache_io_master_M_Cmd),
    .io_master_M_Addr(dcache_io_master_M_Addr),
    .io_master_M_Data(dcache_io_master_M_Data),
    .io_master_M_ByteEn(dcache_io_master_M_ByteEn),
    .io_master_M_AddrSpace(dcache_io_master_M_AddrSpace),
    .io_master_S_Resp(dcache_io_master_S_Resp),
    .io_master_S_Data(dcache_io_master_S_Data),
    .io_slave_M_Cmd(dcache_io_slave_M_Cmd),
    .io_slave_M_Addr(dcache_io_slave_M_Addr),
    .io_slave_M_Data(dcache_io_slave_M_Data),
    .io_slave_M_DataValid(dcache_io_slave_M_DataValid),
    .io_slave_M_DataByteEn(dcache_io_slave_M_DataByteEn),
    .io_slave_S_Resp(dcache_io_slave_S_Resp),
    .io_slave_S_Data(dcache_io_slave_S_Data),
    .io_slave_S_CmdAccept(dcache_io_slave_S_CmdAccept),
    .io_slave_S_DataAccept(dcache_io_slave_S_DataAccept),
    .io_scIO_ena_in(dcache_io_scIO_ena_in),
    .io_scIO_exsc_op(dcache_io_scIO_exsc_op),
    .io_scIO_exsc_opData(dcache_io_scIO_exsc_opData),
    .io_scIO_exsc_opOff(dcache_io_scIO_exsc_opOff),
    .io_scIO_scex_stackTop(dcache_io_scIO_scex_stackTop),
    .io_scIO_scex_memTop(dcache_io_scIO_scex_memTop),
    .io_scIO_illMem(dcache_io_scIO_illMem),
    .io_scIO_stall(dcache_io_scIO_stall),
    .io_invalDCache(dcache_io_invalDCache)
  );
  OcpBurstBus burstBus ( // @[Patmos.scala 107:24]
    .io_master_M_Cmd(burstBus_io_master_M_Cmd),
    .io_master_M_Addr(burstBus_io_master_M_Addr),
    .io_master_M_Data(burstBus_io_master_M_Data),
    .io_master_M_DataValid(burstBus_io_master_M_DataValid),
    .io_master_M_DataByteEn(burstBus_io_master_M_DataByteEn),
    .io_master_S_Resp(burstBus_io_master_S_Resp),
    .io_master_S_Data(burstBus_io_master_S_Data),
    .io_master_S_CmdAccept(burstBus_io_master_S_CmdAccept),
    .io_master_S_DataAccept(burstBus_io_master_S_DataAccept),
    .io_slave_M_Cmd(burstBus_io_slave_M_Cmd),
    .io_slave_M_Addr(burstBus_io_slave_M_Addr),
    .io_slave_M_Data(burstBus_io_slave_M_Data),
    .io_slave_M_DataValid(burstBus_io_slave_M_DataValid),
    .io_slave_M_DataByteEn(burstBus_io_slave_M_DataByteEn),
    .io_slave_S_Resp(burstBus_io_slave_S_Resp),
    .io_slave_S_Data(burstBus_io_slave_S_Data),
    .io_slave_S_CmdAccept(burstBus_io_slave_S_CmdAccept),
    .io_slave_S_DataAccept(burstBus_io_slave_S_DataAccept)
  );
  NoMemoryManagement mmu ( // @[Patmos.scala 119:19]
    .io_virt_M_Cmd(mmu_io_virt_M_Cmd),
    .io_virt_M_Addr(mmu_io_virt_M_Addr),
    .io_virt_M_Data(mmu_io_virt_M_Data),
    .io_virt_M_DataValid(mmu_io_virt_M_DataValid),
    .io_virt_M_DataByteEn(mmu_io_virt_M_DataByteEn),
    .io_virt_S_Resp(mmu_io_virt_S_Resp),
    .io_virt_S_Data(mmu_io_virt_S_Data),
    .io_phys_M_Cmd(mmu_io_phys_M_Cmd),
    .io_phys_M_Addr(mmu_io_phys_M_Addr),
    .io_phys_M_Data(mmu_io_phys_M_Data),
    .io_phys_M_DataValid(mmu_io_phys_M_DataValid),
    .io_phys_M_DataByteEn(mmu_io_phys_M_DataByteEn),
    .io_phys_S_Resp(mmu_io_phys_S_Resp),
    .io_phys_S_Data(mmu_io_phys_S_Data)
  );
  assign io_memPort_M_Cmd = mmu_io_phys_M_Cmd; // @[Patmos.scala 166:14]
  assign io_memPort_M_Addr = mmu_io_phys_M_Addr; // @[Patmos.scala 166:14]
  assign io_memPort_M_Data = mmu_io_phys_M_Data; // @[Patmos.scala 166:14]
  assign io_memPort_M_DataValid = mmu_io_phys_M_DataValid; // @[Patmos.scala 166:14]
  assign io_memPort_M_DataByteEn = mmu_io_phys_M_DataByteEn; // @[Patmos.scala 166:14]
  assign io_memInOut_M_Cmd = memory_io_localInOut_M_Cmd; // @[Patmos.scala 94:15]
  assign io_memInOut_M_Addr = memory_io_localInOut_M_Addr; // @[Patmos.scala 94:15]
  assign io_memInOut_M_Data = memory_io_localInOut_M_Data; // @[Patmos.scala 94:15]
  assign io_memInOut_M_ByteEn = memory_io_localInOut_M_ByteEn; // @[Patmos.scala 94:15]
  assign io_excInOut_S_Resp = exc_io_ocp_S_Resp; // @[Patmos.scala 97:15]
  assign io_excInOut_S_Data = exc_io_ocp_S_Data; // @[Patmos.scala 97:15]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_ena_in = memory_io_ena_out & _T_6; // @[Patmos.scala 127:41]
  assign icache_io_invalidate = exc_io_invalICache; // @[Patmos.scala 148:24]
  assign icache_io_feicache_addrEven = fetch_io_feicache_addrEven; // @[Patmos.scala 66:22]
  assign icache_io_feicache_addrOdd = fetch_io_feicache_addrOdd; // @[Patmos.scala 66:22]
  assign icache_io_exicache_doCallRet = execute_io_exicache_doCallRet; // @[Patmos.scala 68:22]
  assign icache_io_exicache_callRetBase = execute_io_exicache_callRetBase; // @[Patmos.scala 68:22]
  assign icache_io_exicache_callRetAddr = execute_io_exicache_callRetAddr; // @[Patmos.scala 68:22]
  assign icache_io_ocp_port_S_Resp = REG ? 2'h0 : burstBus_io_slave_S_Resp; // @[OcpBurst.scala 159:21 OcpBurst.scala 160:17 OcpBurst.scala 157:10]
  assign icache_io_ocp_port_S_Data = burstBus_io_slave_S_Data; // @[OcpBurst.scala 157:10]
  assign icache_io_ocp_port_S_CmdAccept = burstBus_io_slave_S_CmdAccept; // @[OcpBurst.scala 157:10]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_ena = _T_10 & _T_6; // @[Patmos.scala 131:54]
  assign fetch_io_exfe_doBranch = execute_io_exfe_doBranch; // @[Patmos.scala 88:17]
  assign fetch_io_exfe_branchPc = execute_io_exfe_branchPc; // @[Patmos.scala 88:17]
  assign fetch_io_memfe_doCallRet = memory_io_memfe_doCallRet; // @[Patmos.scala 90:18]
  assign fetch_io_memfe_store = memory_io_memfe_store; // @[Patmos.scala 90:18]
  assign fetch_io_memfe_addr = memory_io_memfe_addr; // @[Patmos.scala 90:18]
  assign fetch_io_memfe_data = memory_io_memfe_data; // @[Patmos.scala 90:18]
  assign fetch_io_icachefe_instrEven = icache_io_icachefe_instrEven; // @[Patmos.scala 67:21]
  assign fetch_io_icachefe_instrOdd = icache_io_icachefe_instrOdd; // @[Patmos.scala 67:21]
  assign fetch_io_icachefe_base = icache_io_icachefe_base; // @[Patmos.scala 67:21]
  assign fetch_io_icachefe_relBase = icache_io_icachefe_relBase; // @[Patmos.scala 67:21]
  assign fetch_io_icachefe_relPc = icache_io_icachefe_relPc; // @[Patmos.scala 67:21]
  assign fetch_io_icachefe_reloc = icache_io_icachefe_reloc; // @[Patmos.scala 67:21]
  assign fetch_io_icachefe_memSel = icache_io_icachefe_memSel; // @[Patmos.scala 67:21]
  assign decode_clock = clock;
  assign decode_reset = reset;
  assign decode_io_ena = _T_10 & _T_6; // @[Patmos.scala 131:54]
  assign decode_io_flush = memory_io_flush | execute_io_brflush; // @[Patmos.scala 144:28]
  assign decode_io_fedec_instr_a = fetch_io_fedec_instr_a; // @[Patmos.scala 71:19]
  assign decode_io_fedec_instr_b = fetch_io_fedec_instr_b; // @[Patmos.scala 71:19]
  assign decode_io_fedec_pc = fetch_io_fedec_pc; // @[Patmos.scala 71:19]
  assign decode_io_fedec_base = fetch_io_fedec_base; // @[Patmos.scala 71:19]
  assign decode_io_fedec_reloc = fetch_io_fedec_reloc; // @[Patmos.scala 71:19]
  assign decode_io_fedec_relPc = fetch_io_fedec_relPc; // @[Patmos.scala 71:19]
  assign decode_io_rfWrite_0_addr = writeback_io_rfWrite_0_addr; // @[Patmos.scala 76:21]
  assign decode_io_rfWrite_0_data = writeback_io_rfWrite_0_data; // @[Patmos.scala 76:21]
  assign decode_io_rfWrite_0_valid = writeback_io_rfWrite_0_valid; // @[Patmos.scala 76:21]
  assign decode_io_rfWrite_1_addr = writeback_io_rfWrite_1_addr; // @[Patmos.scala 76:21]
  assign decode_io_rfWrite_1_data = writeback_io_rfWrite_1_data; // @[Patmos.scala 76:21]
  assign decode_io_rfWrite_1_valid = writeback_io_rfWrite_1_valid; // @[Patmos.scala 76:21]
  assign decode_io_exc_exc = exc_io_excdec_exc; // @[Patmos.scala 99:17]
  assign decode_io_exc_excBase = exc_io_excdec_excBase; // @[Patmos.scala 99:17]
  assign decode_io_exc_excAddr = exc_io_excdec_excAddr; // @[Patmos.scala 99:17]
  assign decode_io_exc_intr = exc_io_excdec_intr; // @[Patmos.scala 99:17]
  assign decode_io_exc_addr = exc_io_excdec_addr; // @[Patmos.scala 99:17]
  assign decode_io_exc_src = exc_io_excdec_src; // @[Patmos.scala 99:17]
  assign decode_io_exc_local = exc_io_excdec_local; // @[Patmos.scala 99:17]
  assign execute_clock = clock;
  assign execute_reset = reset;
  assign execute_io_ena = _T_10 & _T_6; // @[Patmos.scala 131:54]
  assign execute_io_flush = memory_io_flush; // @[Patmos.scala 145:20]
  assign execute_io_decex_base = decode_io_decex_base; // @[Patmos.scala 72:20]
  assign execute_io_decex_relPc = decode_io_decex_relPc; // @[Patmos.scala 72:20]
  assign execute_io_decex_pred_0 = decode_io_decex_pred_0; // @[Patmos.scala 72:20]
  assign execute_io_decex_pred_1 = decode_io_decex_pred_1; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_0_func = decode_io_decex_aluOp_0_func; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_0_isMul = decode_io_decex_aluOp_0_isMul; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_0_isCmp = decode_io_decex_aluOp_0_isCmp; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_0_isPred = decode_io_decex_aluOp_0_isPred; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_0_isBCpy = decode_io_decex_aluOp_0_isBCpy; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_0_isMTS = decode_io_decex_aluOp_0_isMTS; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_0_isMFS = decode_io_decex_aluOp_0_isMFS; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_1_func = decode_io_decex_aluOp_1_func; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_1_isCmp = decode_io_decex_aluOp_1_isCmp; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_1_isPred = decode_io_decex_aluOp_1_isPred; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_1_isBCpy = decode_io_decex_aluOp_1_isBCpy; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_1_isMTS = decode_io_decex_aluOp_1_isMTS; // @[Patmos.scala 72:20]
  assign execute_io_decex_aluOp_1_isMFS = decode_io_decex_aluOp_1_isMFS; // @[Patmos.scala 72:20]
  assign execute_io_decex_predOp_0_func = decode_io_decex_predOp_0_func; // @[Patmos.scala 72:20]
  assign execute_io_decex_predOp_0_dest = decode_io_decex_predOp_0_dest; // @[Patmos.scala 72:20]
  assign execute_io_decex_predOp_0_s1Addr = decode_io_decex_predOp_0_s1Addr; // @[Patmos.scala 72:20]
  assign execute_io_decex_predOp_0_s2Addr = decode_io_decex_predOp_0_s2Addr; // @[Patmos.scala 72:20]
  assign execute_io_decex_predOp_1_func = decode_io_decex_predOp_1_func; // @[Patmos.scala 72:20]
  assign execute_io_decex_predOp_1_dest = decode_io_decex_predOp_1_dest; // @[Patmos.scala 72:20]
  assign execute_io_decex_predOp_1_s1Addr = decode_io_decex_predOp_1_s1Addr; // @[Patmos.scala 72:20]
  assign execute_io_decex_predOp_1_s2Addr = decode_io_decex_predOp_1_s2Addr; // @[Patmos.scala 72:20]
  assign execute_io_decex_jmpOp_branch = decode_io_decex_jmpOp_branch; // @[Patmos.scala 72:20]
  assign execute_io_decex_jmpOp_target = decode_io_decex_jmpOp_target; // @[Patmos.scala 72:20]
  assign execute_io_decex_jmpOp_reloc = decode_io_decex_jmpOp_reloc; // @[Patmos.scala 72:20]
  assign execute_io_decex_memOp_load = decode_io_decex_memOp_load; // @[Patmos.scala 72:20]
  assign execute_io_decex_memOp_store = decode_io_decex_memOp_store; // @[Patmos.scala 72:20]
  assign execute_io_decex_memOp_hword = decode_io_decex_memOp_hword; // @[Patmos.scala 72:20]
  assign execute_io_decex_memOp_byte = decode_io_decex_memOp_byte; // @[Patmos.scala 72:20]
  assign execute_io_decex_memOp_zext = decode_io_decex_memOp_zext; // @[Patmos.scala 72:20]
  assign execute_io_decex_memOp_typ = decode_io_decex_memOp_typ; // @[Patmos.scala 72:20]
  assign execute_io_decex_stackOp = decode_io_decex_stackOp; // @[Patmos.scala 72:20]
  assign execute_io_decex_rsAddr_0 = decode_io_decex_rsAddr_0; // @[Patmos.scala 72:20]
  assign execute_io_decex_rsAddr_1 = decode_io_decex_rsAddr_1; // @[Patmos.scala 72:20]
  assign execute_io_decex_rsAddr_2 = decode_io_decex_rsAddr_2; // @[Patmos.scala 72:20]
  assign execute_io_decex_rsAddr_3 = decode_io_decex_rsAddr_3; // @[Patmos.scala 72:20]
  assign execute_io_decex_rsData_0 = decode_io_decex_rsData_0; // @[Patmos.scala 72:20]
  assign execute_io_decex_rsData_1 = decode_io_decex_rsData_1; // @[Patmos.scala 72:20]
  assign execute_io_decex_rsData_2 = decode_io_decex_rsData_2; // @[Patmos.scala 72:20]
  assign execute_io_decex_rsData_3 = decode_io_decex_rsData_3; // @[Patmos.scala 72:20]
  assign execute_io_decex_rdAddr_0 = decode_io_decex_rdAddr_0; // @[Patmos.scala 72:20]
  assign execute_io_decex_rdAddr_1 = decode_io_decex_rdAddr_1; // @[Patmos.scala 72:20]
  assign execute_io_decex_immVal_0 = decode_io_decex_immVal_0; // @[Patmos.scala 72:20]
  assign execute_io_decex_immVal_1 = decode_io_decex_immVal_1; // @[Patmos.scala 72:20]
  assign execute_io_decex_immOp_0 = decode_io_decex_immOp_0; // @[Patmos.scala 72:20]
  assign execute_io_decex_immOp_1 = decode_io_decex_immOp_1; // @[Patmos.scala 72:20]
  assign execute_io_decex_wrRd_0 = decode_io_decex_wrRd_0; // @[Patmos.scala 72:20]
  assign execute_io_decex_wrRd_1 = decode_io_decex_wrRd_1; // @[Patmos.scala 72:20]
  assign execute_io_decex_callAddr = decode_io_decex_callAddr; // @[Patmos.scala 72:20]
  assign execute_io_decex_call = decode_io_decex_call; // @[Patmos.scala 72:20]
  assign execute_io_decex_ret = decode_io_decex_ret; // @[Patmos.scala 72:20]
  assign execute_io_decex_brcf = decode_io_decex_brcf; // @[Patmos.scala 72:20]
  assign execute_io_decex_trap = decode_io_decex_trap; // @[Patmos.scala 72:20]
  assign execute_io_decex_xcall = decode_io_decex_xcall; // @[Patmos.scala 72:20]
  assign execute_io_decex_xret = decode_io_decex_xret; // @[Patmos.scala 72:20]
  assign execute_io_decex_xsrc = decode_io_decex_xsrc; // @[Patmos.scala 72:20]
  assign execute_io_decex_nonDelayed = decode_io_decex_nonDelayed; // @[Patmos.scala 72:20]
  assign execute_io_decex_illOp = decode_io_decex_illOp; // @[Patmos.scala 72:20]
  assign execute_io_feex_pc = fetch_io_feex_pc; // @[Patmos.scala 92:19]
  assign execute_io_exResult_0_addr = memory_io_exResult_0_addr; // @[Patmos.scala 79:23]
  assign execute_io_exResult_0_data = memory_io_exResult_0_data; // @[Patmos.scala 79:23]
  assign execute_io_exResult_0_valid = memory_io_exResult_0_valid; // @[Patmos.scala 79:23]
  assign execute_io_exResult_1_addr = memory_io_exResult_1_addr; // @[Patmos.scala 79:23]
  assign execute_io_exResult_1_data = memory_io_exResult_1_data; // @[Patmos.scala 79:23]
  assign execute_io_exResult_1_valid = memory_io_exResult_1_valid; // @[Patmos.scala 79:23]
  assign execute_io_memResult_0_addr = writeback_io_memResult_0_addr; // @[Patmos.scala 80:24]
  assign execute_io_memResult_0_data = writeback_io_memResult_0_data; // @[Patmos.scala 80:24]
  assign execute_io_memResult_0_valid = writeback_io_memResult_0_valid; // @[Patmos.scala 80:24]
  assign execute_io_memResult_1_addr = writeback_io_memResult_1_addr; // @[Patmos.scala 80:24]
  assign execute_io_memResult_1_data = writeback_io_memResult_1_data; // @[Patmos.scala 80:24]
  assign execute_io_memResult_1_valid = writeback_io_memResult_1_valid; // @[Patmos.scala 80:24]
  assign execute_io_scex_stackTop = dcache_io_scIO_scex_stackTop; // @[Patmos.scala 84:19]
  assign execute_io_scex_memTop = dcache_io_scIO_scex_memTop; // @[Patmos.scala 84:19]
  assign memory_clock = clock;
  assign memory_reset = reset;
  assign memory_io_ena_in = icache_io_ena_out & ~dcache_io_scIO_stall; // @[Patmos.scala 126:41]
  assign memory_io_exmem_rd_0_addr = execute_io_exmem_rd_0_addr; // @[Patmos.scala 73:19]
  assign memory_io_exmem_rd_0_data = execute_io_exmem_rd_0_data; // @[Patmos.scala 73:19]
  assign memory_io_exmem_rd_0_valid = execute_io_exmem_rd_0_valid; // @[Patmos.scala 73:19]
  assign memory_io_exmem_rd_1_addr = execute_io_exmem_rd_1_addr; // @[Patmos.scala 73:19]
  assign memory_io_exmem_rd_1_data = execute_io_exmem_rd_1_data; // @[Patmos.scala 73:19]
  assign memory_io_exmem_rd_1_valid = execute_io_exmem_rd_1_valid; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_load = execute_io_exmem_mem_load; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_store = execute_io_exmem_mem_store; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_hword = execute_io_exmem_mem_hword; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_byte = execute_io_exmem_mem_byte; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_zext = execute_io_exmem_mem_zext; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_typ = execute_io_exmem_mem_typ; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_addr = execute_io_exmem_mem_addr; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_data = execute_io_exmem_mem_data; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_call = execute_io_exmem_mem_call; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_ret = execute_io_exmem_mem_ret; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_brcf = execute_io_exmem_mem_brcf; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_trap = execute_io_exmem_mem_trap; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_xcall = execute_io_exmem_mem_xcall; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_xret = execute_io_exmem_mem_xret; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_xsrc = execute_io_exmem_mem_xsrc; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_illOp = execute_io_exmem_mem_illOp; // @[Patmos.scala 73:19]
  assign memory_io_exmem_mem_nonDelayed = execute_io_exmem_mem_nonDelayed; // @[Patmos.scala 73:19]
  assign memory_io_exmem_base = execute_io_exmem_base; // @[Patmos.scala 73:19]
  assign memory_io_exmem_relPc = execute_io_exmem_relPc; // @[Patmos.scala 73:19]
  assign memory_io_localInOut_S_Resp = io_memInOut_S_Resp; // @[Patmos.scala 94:15]
  assign memory_io_localInOut_S_Data = io_memInOut_S_Data; // @[Patmos.scala 94:15]
  assign memory_io_globalInOut_S_Resp = dcache_io_master_S_Resp; // @[Patmos.scala 104:27]
  assign memory_io_globalInOut_S_Data = dcache_io_master_S_Data; // @[Patmos.scala 104:27]
  assign memory_io_icacheIllMem = icache_io_illMem; // @[Patmos.scala 69:26]
  assign memory_io_scacheIllMem = dcache_io_scIO_illMem; // @[Patmos.scala 85:26]
  assign writeback_io_memwb_rd_0_addr = memory_io_memwb_rd_0_addr; // @[Patmos.scala 74:22]
  assign writeback_io_memwb_rd_0_data = memory_io_memwb_rd_0_data; // @[Patmos.scala 74:22]
  assign writeback_io_memwb_rd_0_valid = memory_io_memwb_rd_0_valid; // @[Patmos.scala 74:22]
  assign writeback_io_memwb_rd_1_addr = memory_io_memwb_rd_1_addr; // @[Patmos.scala 74:22]
  assign writeback_io_memwb_rd_1_data = memory_io_memwb_rd_1_data; // @[Patmos.scala 74:22]
  assign writeback_io_memwb_rd_1_valid = memory_io_memwb_rd_1_valid; // @[Patmos.scala 74:22]
  assign exc_clock = clock;
  assign exc_reset = reset;
  assign exc_io_ena = _T_10 & _T_6; // @[Patmos.scala 131:54]
  assign exc_io_ocp_M_Cmd = io_excInOut_M_Cmd; // @[Patmos.scala 97:15]
  assign exc_io_ocp_M_Addr = io_excInOut_M_Addr; // @[Patmos.scala 97:15]
  assign exc_io_ocp_M_Data = io_excInOut_M_Data; // @[Patmos.scala 97:15]
  assign exc_io_intrs_0 = io_interrupts_0; // @[Patmos.scala 98:16]
  assign exc_io_intrs_1 = io_interrupts_1; // @[Patmos.scala 98:16]
  assign exc_io_intrs_2 = io_interrupts_2; // @[Patmos.scala 98:16]
  assign exc_io_intrs_3 = io_interrupts_3; // @[Patmos.scala 98:16]
  assign exc_io_intrs_4 = io_interrupts_4; // @[Patmos.scala 98:16]
  assign exc_io_intrs_5 = io_interrupts_5; // @[Patmos.scala 98:16]
  assign exc_io_memexc_call = memory_io_exc_call; // @[Patmos.scala 100:17]
  assign exc_io_memexc_ret = memory_io_exc_ret; // @[Patmos.scala 100:17]
  assign exc_io_memexc_src = memory_io_exc_src; // @[Patmos.scala 100:17]
  assign exc_io_memexc_exc = memory_io_exc_exc; // @[Patmos.scala 100:17]
  assign exc_io_memexc_excBase = memory_io_exc_excBase; // @[Patmos.scala 100:17]
  assign exc_io_memexc_excAddr = memory_io_exc_excAddr; // @[Patmos.scala 100:17]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_master_M_Cmd = memory_io_globalInOut_M_Cmd; // @[Patmos.scala 103:22]
  assign dcache_io_master_M_Addr = memory_io_globalInOut_M_Addr; // @[Patmos.scala 103:22]
  assign dcache_io_master_M_Data = memory_io_globalInOut_M_Data; // @[Patmos.scala 103:22]
  assign dcache_io_master_M_ByteEn = memory_io_globalInOut_M_ByteEn; // @[Patmos.scala 103:22]
  assign dcache_io_master_M_AddrSpace = memory_io_globalInOut_M_AddrSpace; // @[Patmos.scala 103:22]
  assign dcache_io_slave_S_Resp = REG ? burstBus_io_slave_S_Resp : 2'h0; // @[OcpBurst.scala 159:21 OcpBurst.scala 156:11 OcpBurst.scala 163:18]
  assign dcache_io_slave_S_Data = burstBus_io_slave_S_Data; // @[OcpBurst.scala 156:11]
  assign dcache_io_slave_S_CmdAccept = burstBus_io_slave_S_CmdAccept; // @[OcpBurst.scala 156:11]
  assign dcache_io_slave_S_DataAccept = burstBus_io_slave_S_DataAccept; // @[OcpBurst.scala 156:11]
  assign dcache_io_scIO_ena_in = memory_io_ena_out & icache_io_ena_out; // @[Patmos.scala 128:46]
  assign dcache_io_scIO_exsc_op = execute_io_exsc_op; // @[Patmos.scala 83:23]
  assign dcache_io_scIO_exsc_opData = execute_io_exsc_opData; // @[Patmos.scala 83:23]
  assign dcache_io_scIO_exsc_opOff = execute_io_exsc_opOff; // @[Patmos.scala 83:23]
  assign dcache_io_invalDCache = exc_io_invalDCache; // @[Patmos.scala 149:25]
  assign burstBus_io_master_S_Resp = mmu_io_virt_S_Resp; // @[Patmos.scala 123:24]
  assign burstBus_io_master_S_Data = mmu_io_virt_S_Data; // @[Patmos.scala 123:24]
  assign burstBus_io_master_S_CmdAccept = 1'h1; // @[Patmos.scala 123:24]
  assign burstBus_io_master_S_DataAccept = 1'h1; // @[Patmos.scala 123:24]
  assign burstBus_io_slave_M_Cmd = dcache_io_slave_M_Cmd | icache_io_ocp_port_M_Cmd; // @[OcpBurst.scala 154:31]
  assign burstBus_io_slave_M_Addr = _T_3 ? dcache_io_slave_M_Addr : icache_io_ocp_port_M_Addr; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign burstBus_io_slave_M_Data = _T_3 ? dcache_io_slave_M_Data : 32'h0; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign burstBus_io_slave_M_DataValid = _T_3 & dcache_io_slave_M_DataValid; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign burstBus_io_slave_M_DataByteEn = _T_3 ? dcache_io_slave_M_DataByteEn : 4'hf; // @[OcpBurst.scala 151:19 OcpBurst.scala 152:14 OcpBurst.scala 150:12]
  assign mmu_io_virt_M_Cmd = burstBus_io_master_M_Cmd; // @[Patmos.scala 122:17]
  assign mmu_io_virt_M_Addr = burstBus_io_master_M_Addr; // @[Patmos.scala 122:17]
  assign mmu_io_virt_M_Data = burstBus_io_master_M_Data; // @[Patmos.scala 122:17]
  assign mmu_io_virt_M_DataValid = burstBus_io_master_M_DataValid; // @[Patmos.scala 122:17]
  assign mmu_io_virt_M_DataByteEn = burstBus_io_master_M_DataByteEn; // @[Patmos.scala 122:17]
  assign mmu_io_phys_S_Resp = io_memPort_S_Resp; // @[Patmos.scala 166:14]
  assign mmu_io_phys_S_Data = io_memPort_S_Data; // @[Patmos.scala 166:14]
  always @(posedge clock) begin
    if (icache_io_ocp_port_M_Cmd != 3'h0) begin // @[OcpBurst.scala 146:18]
      REG <= 1'h0;
    end else begin
      REG <= _T_2;
    end
    enableReg <= _T_10 & _T_6; // @[Patmos.scala 131:54]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  enableReg = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HardlockOCPWrapper(
  input        clock,
  input        reset,
  input  [2:0] io_cores_0_M_Cmd,
  output [1:0] io_cores_0_S_Resp
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  reqReg; // @[Hardlock.scala 84:19]
  wire  _GEN_1 = reqReg ? 1'h0 : reqReg; // @[Hardlock.scala 101:86 Hardlock.scala 102:19 Hardlock.scala 87:12]
  wire  reqBools_0 = io_cores_0_M_Cmd != 3'h0 | _GEN_1; // @[Hardlock.scala 97:45 Hardlock.scala 98:19]
  assign io_cores_0_S_Resp = reqReg ? 2'h1 : 2'h0; // @[Hardlock.scala 107:81 Hardlock.scala 108:26 Hardlock.scala 106:24]
  always @(posedge clock) begin
    if (reset) begin // @[Hardlock.scala 84:19]
      reqReg <= 1'h0; // @[Hardlock.scala 84:19]
    end else if (io_cores_0_M_Cmd != 3'h0) begin // @[Hardlock.scala 97:45]
      reqReg <= reqBools_0; // @[Hardlock.scala 99:14]
    end else if (reqReg) begin // @[Hardlock.scala 101:86]
      reqReg <= reqBools_0; // @[Hardlock.scala 103:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reqReg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module QueueCompatibility(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:15]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Uart(
  input         clock,
  input         reset,
  input  [2:0]  io_ocp_M_Cmd,
  input  [31:0] io_ocp_M_Addr,
  input  [31:0] io_ocp_M_Data,
  output [1:0]  io_ocp_S_Resp,
  output [31:0] io_ocp_S_Data,
  output        io_pins_tx,
  input         io_pins_rx
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  txQueue_clock; // @[Uart.scala 58:25]
  wire  txQueue_reset; // @[Uart.scala 58:25]
  wire  txQueue_io_enq_ready; // @[Uart.scala 58:25]
  wire  txQueue_io_enq_valid; // @[Uart.scala 58:25]
  wire [7:0] txQueue_io_enq_bits; // @[Uart.scala 58:25]
  wire  txQueue_io_deq_ready; // @[Uart.scala 58:25]
  wire  txQueue_io_deq_valid; // @[Uart.scala 58:25]
  wire [7:0] txQueue_io_deq_bits; // @[Uart.scala 58:25]
  wire  rxQueue_clock; // @[Uart.scala 76:25]
  wire  rxQueue_reset; // @[Uart.scala 76:25]
  wire  rxQueue_io_enq_ready; // @[Uart.scala 76:25]
  wire  rxQueue_io_enq_valid; // @[Uart.scala 76:25]
  wire [7:0] rxQueue_io_enq_bits; // @[Uart.scala 76:25]
  wire  rxQueue_io_deq_ready; // @[Uart.scala 76:25]
  wire  rxQueue_io_deq_valid; // @[Uart.scala 76:25]
  wire [7:0] rxQueue_io_deq_bits; // @[Uart.scala 76:25]
  reg [9:0] tx_baud_counter; // @[Uart.scala 49:34]
  reg  tx_baud_tick; // @[Uart.scala 50:34]
  reg  tx_state; // @[Uart.scala 53:34]
  reg [9:0] tx_buff; // @[Uart.scala 54:34]
  reg  tx_reg; // @[Uart.scala 55:34]
  reg [3:0] tx_counter; // @[Uart.scala 56:34]
  reg  rxd_reg0; // @[Uart.scala 63:34]
  reg  rxd_reg1; // @[Uart.scala 64:34]
  reg  rxd_reg2; // @[Uart.scala 65:34]
  reg [9:0] rx_baud_counter; // @[Uart.scala 67:34]
  reg  rx_baud_tick; // @[Uart.scala 68:34]
  reg  rx_enable; // @[Uart.scala 69:34]
  reg [7:0] rx_buff; // @[Uart.scala 71:34]
  reg [2:0] rx_counter; // @[Uart.scala 72:34]
  reg [1:0] rx_state; // @[Uart.scala 74:34]
  reg [1:0] respReg; // @[Uart.scala 82:22]
  reg [7:0] rdDataReg; // @[Uart.scala 85:24]
  wire [7:0] _T_3 = {6'h0,rxQueue_io_deq_valid,txQueue_io_enq_ready}; // @[Cat.scala 30:58]
  wire  _T_10 = tx_baud_counter == 10'h2b6; // @[Uart.scala 108:27]
  wire [9:0] _T_12 = tx_baud_counter + 10'h1; // @[Uart.scala 113:48]
  wire [8:0] hi_1 = {1'h1,txQueue_io_deq_bits}; // @[Cat.scala 30:58]
  wire [9:0] _T_14 = {1'h1,txQueue_io_deq_bits,1'h0}; // @[Cat.scala 30:58]
  wire  _GEN_7 = txQueue_io_deq_valid; // @[Uart.scala 120:37 Uart.scala 121:32 Uart.scala 61:29]
  wire [9:0] _GEN_8 = txQueue_io_deq_valid ? _T_14 : tx_buff; // @[Uart.scala 120:37 Uart.scala 122:32 Uart.scala 54:34]
  wire  _GEN_9 = txQueue_io_deq_valid | tx_state; // @[Uart.scala 120:37 Uart.scala 123:32 Uart.scala 53:34]
  wire  _GEN_10 = ~tx_state & _GEN_7; // @[Uart.scala 119:33 Uart.scala 61:29]
  wire [9:0] _GEN_11 = ~tx_state ? _GEN_8 : tx_buff; // @[Uart.scala 119:33 Uart.scala 54:34]
  wire  _GEN_12 = ~tx_state ? _GEN_9 : tx_state; // @[Uart.scala 119:33 Uart.scala 53:34]
  wire [8:0] lo = tx_buff[9:1]; // @[Uart.scala 129:54]
  wire [9:0] _T_17 = {1'h0,lo}; // @[Cat.scala 30:58]
  wire  _T_19 = tx_counter == 4'ha; // @[Uart.scala 131:47]
  wire [3:0] _T_21 = tx_counter + 4'h1; // @[Uart.scala 131:81]
  wire [3:0] _T_22 = tx_counter == 4'ha ? 4'h0 : _T_21; // @[Uart.scala 131:35]
  wire  _GEN_13 = txQueue_io_deq_valid | _GEN_10; // @[Uart.scala 134:43 Uart.scala 135:38]
  wire [9:0] _GEN_14 = txQueue_io_deq_valid ? {{1'd0}, hi_1} : _T_17; // @[Uart.scala 134:43 Uart.scala 136:38 Uart.scala 129:29]
  wire  _GEN_15 = txQueue_io_deq_valid ? 1'h0 : 1'h1; // @[Uart.scala 134:43 Uart.scala 137:38 Uart.scala 141:33]
  wire  _GEN_16 = txQueue_io_deq_valid & _GEN_12; // @[Uart.scala 134:43 Uart.scala 143:33]
  wire  _GEN_17 = _T_19 ? _GEN_13 : _GEN_10; // @[Uart.scala 133:44]
  wire  _GEN_19 = _T_19 ? _GEN_15 : tx_buff[0]; // @[Uart.scala 133:44 Uart.scala 130:29]
  wire  _GEN_23 = tx_baud_tick ? _GEN_19 : tx_reg; // @[Uart.scala 128:40 Uart.scala 55:34]
  wire  _GEN_25 = tx_baud_tick ? _GEN_17 : _GEN_10; // @[Uart.scala 128:40]
  wire  _GEN_28 = tx_state ? _GEN_23 : tx_reg; // @[Uart.scala 127:33 Uart.scala 55:34]
  wire  _T_25 = rx_baud_counter == 10'h2b6; // @[Uart.scala 155:31]
  wire [9:0] _T_27 = rx_baud_counter + 10'h1; // @[Uart.scala 160:52]
  wire [9:0] _GEN_32 = rx_baud_counter == 10'h2b6 ? 10'h0 : _T_27; // @[Uart.scala 155:60 Uart.scala 156:33 Uart.scala 160:33]
  wire [9:0] _GEN_34 = rx_enable ? _GEN_32 : rx_baud_counter; // @[Uart.scala 154:22 Uart.scala 67:34]
  wire  _T_29 = ~rxd_reg2; // @[Uart.scala 175:24]
  wire [9:0] _T_30 = 10'h2b6 / 10'h2; // @[Uart.scala 177:57]
  wire [1:0] _GEN_36 = ~rxd_reg2 ? 2'h1 : rx_state; // @[Uart.scala 175:36 Uart.scala 176:29 Uart.scala 74:34]
  wire  _GEN_38 = ~rxd_reg2 | rx_enable; // @[Uart.scala 175:36 Uart.scala 178:29 Uart.scala 69:34]
  wire [1:0] _GEN_39 = rx_state == 2'h0 ? _GEN_36 : rx_state; // @[Uart.scala 174:33 Uart.scala 74:34]
  wire  _GEN_41 = rx_state == 2'h0 ? _GEN_38 : rx_enable; // @[Uart.scala 174:33 Uart.scala 69:34]
  wire [1:0] _GEN_42 = _T_29 ? 2'h2 : 2'h0; // @[Uart.scala 184:41 Uart.scala 185:33 Uart.scala 188:33]
  wire [1:0] _GEN_43 = rx_baud_tick ? _GEN_42 : _GEN_39; // @[Uart.scala 183:41]
  wire [1:0] _GEN_44 = rx_state == 2'h1 ? _GEN_43 : _GEN_39; // @[Uart.scala 182:33]
  wire  _T_36 = rx_counter == 3'h7; // @[Uart.scala 195:40]
  wire [1:0] _T_37 = rx_counter == 3'h7 ? 2'h3 : 2'h2; // @[Uart.scala 195:28]
  wire [2:0] _T_40 = rx_counter + 3'h1; // @[Uart.scala 196:75]
  wire [6:0] lo_1 = rx_buff[7:1]; // @[Uart.scala 197:46]
  wire [7:0] _T_42 = {rxd_reg2,lo_1}; // @[Cat.scala 30:58]
  wire [1:0] _GEN_45 = rx_baud_tick ? _T_37 : _GEN_44; // @[Uart.scala 194:40 Uart.scala 195:22]
  wire [1:0] _GEN_48 = rx_state == 2'h2 ? _GEN_45 : _GEN_44; // @[Uart.scala 193:41]
  wire  _GEN_58 = rx_baud_tick & rxd_reg2; // @[Uart.scala 202:40 Uart.scala 78:29]
  wire [2:0] uartOcpEmu_Cmd = io_ocp_M_Cmd; // @[Uart.scala 44:26 Uart.scala 46:16]
  wire [31:0] uartOcpEmu_Addr = io_ocp_M_Addr; // @[Uart.scala 44:26 Uart.scala 46:16]
  wire [31:0] uartOcpEmu_Data = io_ocp_M_Data; // @[Uart.scala 44:26 Uart.scala 46:16]
  QueueCompatibility txQueue ( // @[Uart.scala 58:25]
    .clock(txQueue_clock),
    .reset(txQueue_reset),
    .io_enq_ready(txQueue_io_enq_ready),
    .io_enq_valid(txQueue_io_enq_valid),
    .io_enq_bits(txQueue_io_enq_bits),
    .io_deq_ready(txQueue_io_deq_ready),
    .io_deq_valid(txQueue_io_deq_valid),
    .io_deq_bits(txQueue_io_deq_bits)
  );
  QueueCompatibility rxQueue ( // @[Uart.scala 76:25]
    .clock(rxQueue_clock),
    .reset(rxQueue_reset),
    .io_enq_ready(rxQueue_io_enq_ready),
    .io_enq_valid(rxQueue_io_enq_valid),
    .io_enq_bits(rxQueue_io_enq_bits),
    .io_deq_ready(rxQueue_io_deq_ready),
    .io_deq_valid(rxQueue_io_deq_valid),
    .io_deq_bits(rxQueue_io_deq_bits)
  );
  assign io_ocp_S_Resp = respReg; // @[Uart.scala 104:19]
  assign io_ocp_S_Data = {{24'd0}, rdDataReg}; // @[Uart.scala 105:19]
  assign io_pins_tx = tx_reg; // @[Uart.scala 150:16]
  assign txQueue_clock = clock;
  assign txQueue_reset = reset;
  assign txQueue_io_enq_valid = io_ocp_M_Cmd == 3'h1; // @[Uart.scala 91:24]
  assign txQueue_io_enq_bits = io_ocp_M_Cmd == 3'h1 ? io_ocp_M_Data[7:0] : io_ocp_M_Data[7:0]; // @[Uart.scala 91:39 Uart.scala 93:29 Uart.scala 59:29]
  assign txQueue_io_deq_ready = tx_state ? _GEN_25 : _GEN_10; // @[Uart.scala 127:33]
  assign rxQueue_clock = clock;
  assign rxQueue_reset = reset;
  assign rxQueue_io_enq_valid = rx_state == 2'h3 & _GEN_58; // @[Uart.scala 201:37 Uart.scala 78:29]
  assign rxQueue_io_enq_bits = rx_buff; // @[Uart.scala 201:37 Uart.scala 77:29]
  assign rxQueue_io_deq_ready = io_ocp_M_Cmd == 3'h2 & io_ocp_M_Addr[2]; // @[Uart.scala 98:38 Uart.scala 100:30 Uart.scala 79:29]
  always @(posedge clock) begin
    if (reset) begin // @[Uart.scala 49:34]
      tx_baud_counter <= 10'h0; // @[Uart.scala 49:34]
    end else if (tx_baud_counter == 10'h2b6) begin // @[Uart.scala 108:56]
      tx_baud_counter <= 10'h0; // @[Uart.scala 109:29]
    end else begin
      tx_baud_counter <= _T_12; // @[Uart.scala 113:29]
    end
    if (reset) begin // @[Uart.scala 50:34]
      tx_baud_tick <= 1'h0; // @[Uart.scala 50:34]
    end else begin
      tx_baud_tick <= _T_10;
    end
    if (reset) begin // @[Uart.scala 53:34]
      tx_state <= 1'h0; // @[Uart.scala 53:34]
    end else if (tx_state) begin // @[Uart.scala 127:33]
      if (tx_baud_tick) begin // @[Uart.scala 128:40]
        if (_T_19) begin // @[Uart.scala 133:44]
          tx_state <= _GEN_16;
        end else begin
          tx_state <= _GEN_12;
        end
      end else begin
        tx_state <= _GEN_12;
      end
    end else begin
      tx_state <= _GEN_12;
    end
    if (reset) begin // @[Uart.scala 54:34]
      tx_buff <= 10'h0; // @[Uart.scala 54:34]
    end else if (tx_state) begin // @[Uart.scala 127:33]
      if (tx_baud_tick) begin // @[Uart.scala 128:40]
        if (_T_19) begin // @[Uart.scala 133:44]
          tx_buff <= _GEN_14;
        end else begin
          tx_buff <= _T_17; // @[Uart.scala 129:29]
        end
      end else begin
        tx_buff <= _GEN_11;
      end
    end else begin
      tx_buff <= _GEN_11;
    end
    tx_reg <= reset | _GEN_28; // @[Uart.scala 55:34 Uart.scala 55:34]
    if (reset) begin // @[Uart.scala 56:34]
      tx_counter <= 4'h0; // @[Uart.scala 56:34]
    end else if (tx_state) begin // @[Uart.scala 127:33]
      if (tx_baud_tick) begin // @[Uart.scala 128:40]
        if (tx_counter == 4'ha) begin // @[Uart.scala 133:44]
          tx_counter <= {{3'd0}, _GEN_7};
        end else begin
          tx_counter <= _T_22; // @[Uart.scala 131:29]
        end
      end
    end
    rxd_reg0 <= reset | io_pins_rx; // @[Uart.scala 63:34 Uart.scala 63:34 Uart.scala 168:29]
    rxd_reg1 <= reset | rxd_reg0; // @[Uart.scala 64:34 Uart.scala 64:34 Uart.scala 169:29]
    rxd_reg2 <= reset | rxd_reg1; // @[Uart.scala 65:34 Uart.scala 65:34 Uart.scala 170:29]
    if (reset) begin // @[Uart.scala 67:34]
      rx_baud_counter <= 10'h0; // @[Uart.scala 67:34]
    end else if (rx_state == 2'h0) begin // @[Uart.scala 174:33]
      if (~rxd_reg2) begin // @[Uart.scala 175:36]
        rx_baud_counter <= _T_30; // @[Uart.scala 177:29]
      end else begin
        rx_baud_counter <= _GEN_34;
      end
    end else begin
      rx_baud_counter <= _GEN_34;
    end
    if (reset) begin // @[Uart.scala 68:34]
      rx_baud_tick <= 1'h0; // @[Uart.scala 68:34]
    end else if (rx_enable) begin // @[Uart.scala 154:22]
      rx_baud_tick <= _T_25;
    end
    if (reset) begin // @[Uart.scala 69:34]
      rx_enable <= 1'h0; // @[Uart.scala 69:34]
    end else if (rx_state == 2'h3) begin // @[Uart.scala 201:37]
      if (rx_baud_tick) begin // @[Uart.scala 202:40]
        rx_enable <= 1'h0;
      end else begin
        rx_enable <= _GEN_41;
      end
    end else begin
      rx_enable <= _GEN_41;
    end
    if (reset) begin // @[Uart.scala 71:34]
      rx_buff <= 8'h0; // @[Uart.scala 71:34]
    end else if (rx_state == 2'h2) begin // @[Uart.scala 193:41]
      if (rx_baud_tick) begin // @[Uart.scala 194:40]
        rx_buff <= _T_42; // @[Uart.scala 197:21]
      end
    end
    if (reset) begin // @[Uart.scala 72:34]
      rx_counter <= 3'h0; // @[Uart.scala 72:34]
    end else if (rx_state == 2'h2) begin // @[Uart.scala 193:41]
      if (rx_baud_tick) begin // @[Uart.scala 194:40]
        if (_T_36) begin // @[Uart.scala 196:30]
          rx_counter <= 3'h0;
        end else begin
          rx_counter <= _T_40;
        end
      end
    end
    if (reset) begin // @[Uart.scala 74:34]
      rx_state <= 2'h0; // @[Uart.scala 74:34]
    end else if (rx_state == 2'h3) begin // @[Uart.scala 201:37]
      if (rx_baud_tick) begin // @[Uart.scala 202:40]
        rx_state <= 2'h0;
      end else begin
        rx_state <= _GEN_48;
      end
    end else begin
      rx_state <= _GEN_48;
    end
    if (reset) begin // @[Uart.scala 82:22]
      respReg <= 2'h0; // @[Uart.scala 82:22]
    end else if (io_ocp_M_Cmd == 3'h2) begin // @[Uart.scala 98:38]
      respReg <= 2'h1; // @[Uart.scala 99:17]
    end else if (io_ocp_M_Cmd == 3'h1) begin // @[Uart.scala 91:39]
      respReg <= 2'h1; // @[Uart.scala 92:17]
    end else begin
      respReg <= 2'h0; // @[Uart.scala 83:13]
    end
    if (reset) begin // @[Uart.scala 85:24]
      rdDataReg <= 8'h0; // @[Uart.scala 85:24]
    end else if (~io_ocp_M_Addr[2]) begin // @[Uart.scala 86:21]
      rdDataReg <= _T_3;
    end else begin
      rdDataReg <= rxQueue_io_deq_bits;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tx_baud_counter = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  tx_baud_tick = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  tx_state = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  tx_buff = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  tx_reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  tx_counter = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  rxd_reg0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  rxd_reg1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  rxd_reg2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  rx_baud_counter = _RAND_9[9:0];
  _RAND_10 = {1{`RANDOM}};
  rx_baud_tick = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  rx_enable = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  rx_buff = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  rx_counter = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  rx_state = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  respReg = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  rdDataReg = _RAND_16[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module UartCmp(
  input         clock,
  input         reset,
  input  [2:0]  io_cores_0_M_Cmd,
  input  [31:0] io_cores_0_M_Addr,
  input  [31:0] io_cores_0_M_Data,
  output [1:0]  io_cores_0_S_Resp,
  output [31:0] io_cores_0_S_Data,
  output        io_pins_tx,
  input         io_pins_rx
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  uart_clock; // @[UartCmp.scala 29:20]
  wire  uart_reset; // @[UartCmp.scala 29:20]
  wire [2:0] uart_io_ocp_M_Cmd; // @[UartCmp.scala 29:20]
  wire [31:0] uart_io_ocp_M_Addr; // @[UartCmp.scala 29:20]
  wire [31:0] uart_io_ocp_M_Data; // @[UartCmp.scala 29:20]
  wire [1:0] uart_io_ocp_S_Resp; // @[UartCmp.scala 29:20]
  wire [31:0] uart_io_ocp_S_Data; // @[UartCmp.scala 29:20]
  wire  uart_io_pins_tx; // @[UartCmp.scala 29:20]
  wire  uart_io_pins_rx; // @[UartCmp.scala 29:20]
  wire  _T = io_cores_0_M_Cmd != 3'h0; // @[UartCmp.scala 33:59]
  reg  REG; // @[UartCmp.scala 36:21]
  wire  _GEN_0 = uart_io_ocp_S_Resp == 2'h1 ? 1'h0 : REG; // @[UartCmp.scala 39:52 UartCmp.scala 40:14 UartCmp.scala 36:21]
  wire  _GEN_1 = _T | _GEN_0; // @[UartCmp.scala 37:45 UartCmp.scala 38:14]
  Uart uart ( // @[UartCmp.scala 29:20]
    .clock(uart_clock),
    .reset(uart_reset),
    .io_ocp_M_Cmd(uart_io_ocp_M_Cmd),
    .io_ocp_M_Addr(uart_io_ocp_M_Addr),
    .io_ocp_M_Data(uart_io_ocp_M_Data),
    .io_ocp_S_Resp(uart_io_ocp_S_Resp),
    .io_ocp_S_Data(uart_io_ocp_S_Data),
    .io_pins_tx(uart_io_pins_tx),
    .io_pins_rx(uart_io_pins_rx)
  );
  assign io_cores_0_S_Resp = ~REG ? 2'h0 : uart_io_ocp_S_Resp; // @[UartCmp.scala 45:33 UartCmp.scala 46:26 UartCmp.scala 44:24]
  assign io_cores_0_S_Data = uart_io_ocp_S_Data; // @[UartCmp.scala 43:24]
  assign io_pins_tx = uart_io_pins_tx; // @[UartCmp.scala 31:11]
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_io_ocp_M_Cmd = io_cores_0_M_Cmd; // @[UartCmp.scala 33:17]
  assign uart_io_ocp_M_Addr = io_cores_0_M_Addr; // @[UartCmp.scala 33:17]
  assign uart_io_ocp_M_Data = io_cores_0_M_Data; // @[UartCmp.scala 33:17]
  assign uart_io_pins_rx = io_pins_rx; // @[UartCmp.scala 31:11]
  always @(posedge clock) begin
    if (reset) begin // @[UartCmp.scala 36:21]
      REG <= 1'h0; // @[UartCmp.scala 36:21]
    end else begin
      REG <= _GEN_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CpuInfo(
  input         clock,
  input  [2:0]  io_ocp_M_Cmd,
  input  [31:0] io_ocp_M_Addr,
  output [1:0]  io_ocp_S_Resp,
  output [31:0] io_ocp_S_Data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] masterReg_Cmd; // @[CpuInfo.scala 26:22]
  reg [31:0] masterReg_Addr; // @[CpuInfo.scala 26:22]
  wire [1:0] _GEN_0 = masterReg_Cmd == 3'h1 ? 2'h1 : 2'h0; // @[CpuInfo.scala 35:37 CpuInfo.scala 36:10 CpuInfo.scala 31:8]
  wire  _T_3 = 4'h0 == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_4 = 4'h1 == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_5 = 4'h2 == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_6 = 4'h3 == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_7 = 4'h4 == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_8 = 4'h5 == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_11 = 4'h6 == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_12 = 4'h7 == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_15 = 4'h8 == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_16 = 4'h9 == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_20 = 4'ha == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_21 = 4'hb == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_22 = 4'hc == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire  _T_23 = 4'hd == masterReg_Addr[5:2]; // @[Conditional.scala 37:30]
  wire [11:0] _GEN_1 = _T_23 ? 12'h800 : 12'h0; // @[Conditional.scala 39:67 CpuInfo.scala 74:30 CpuInfo.scala 32:8]
  wire [11:0] _GEN_2 = _T_22 ? 12'h400 : _GEN_1; // @[Conditional.scala 39:67 CpuInfo.scala 71:30]
  wire [11:0] _GEN_3 = _T_21 ? 12'h0 : _GEN_2; // @[Conditional.scala 39:67 CpuInfo.scala 68:30]
  wire [11:0] _GEN_4 = _T_20 ? 12'h800 : _GEN_3; // @[Conditional.scala 39:67 CpuInfo.scala 66:30]
  wire [31:0] _GEN_5 = _T_16 ? 32'h1000001 : {{20'd0}, _GEN_4}; // @[Conditional.scala 39:67 CpuInfo.scala 63:30]
  wire [31:0] _GEN_6 = _T_15 ? 32'h1000 : _GEN_5; // @[Conditional.scala 39:67 CpuInfo.scala 61:30]
  wire [31:0] _GEN_7 = _T_12 ? 32'h1020010 : _GEN_6; // @[Conditional.scala 39:67 CpuInfo.scala 58:30]
  wire [31:0] _GEN_8 = _T_11 ? 32'h2000 : _GEN_7; // @[Conditional.scala 39:67 CpuInfo.scala 56:30]
  wire [31:0] _GEN_9 = _T_8 ? 32'h400 : _GEN_8; // @[Conditional.scala 39:67 CpuInfo.scala 53:30]
  wire [31:0] _GEN_10 = _T_7 ? 32'h200000 : _GEN_9; // @[Conditional.scala 39:67 CpuInfo.scala 51:30]
  wire [31:0] _GEN_11 = _T_6 ? 32'h2 : _GEN_10; // @[Conditional.scala 39:67 CpuInfo.scala 48:30]
  wire [31:0] _GEN_12 = _T_5 ? 32'h1 : _GEN_11; // @[Conditional.scala 39:67 CpuInfo.scala 47:30]
  wire [31:0] _GEN_13 = _T_4 ? 32'h4c4b400 : _GEN_12; // @[Conditional.scala 39:67 CpuInfo.scala 46:30]
  wire [31:0] _GEN_14 = _T_3 ? 32'h0 : _GEN_13; // @[Conditional.scala 40:58 CpuInfo.scala 45:30]
  wire [31:0] _GEN_16 = 4'h1 == masterReg_Addr[5:2] ? 32'h0 : 32'hf0008024; // @[CpuInfo.scala 77:10 CpuInfo.scala 77:10]
  wire [31:0] _GEN_17 = 4'h2 == masterReg_Addr[5:2] ? 32'h20000 : _GEN_16; // @[CpuInfo.scala 77:10 CpuInfo.scala 77:10]
  wire [31:0] _GEN_18 = 4'h3 == masterReg_Addr[5:2] ? 32'h40c : _GEN_17; // @[CpuInfo.scala 77:10 CpuInfo.scala 77:10]
  wire [31:0] _GEN_19 = 4'h4 == masterReg_Addr[5:2] ? 32'h70c : _GEN_18; // @[CpuInfo.scala 77:10 CpuInfo.scala 77:10]
  wire [31:0] _GEN_20 = 4'h5 == masterReg_Addr[5:2] ? 32'h6bc : _GEN_19; // @[CpuInfo.scala 77:10 CpuInfo.scala 77:10]
  wire [31:0] _GEN_21 = 4'h6 == masterReg_Addr[5:2] ? 32'h6f0 : _GEN_20; // @[CpuInfo.scala 77:10 CpuInfo.scala 77:10]
  wire [31:0] _GEN_22 = 4'h7 == masterReg_Addr[5:2] ? 32'h6f8 : _GEN_21; // @[CpuInfo.scala 77:10 CpuInfo.scala 77:10]
  wire [31:0] _GEN_23 = 4'h8 == masterReg_Addr[5:2] ? 32'h700 : _GEN_22; // @[CpuInfo.scala 77:10 CpuInfo.scala 77:10]
  assign io_ocp_S_Resp = masterReg_Cmd == 3'h2 ? 2'h1 : _GEN_0; // @[CpuInfo.scala 80:37 CpuInfo.scala 81:10]
  assign io_ocp_S_Data = masterReg_Addr[15] ? _GEN_23 : _GEN_14; // @[CpuInfo.scala 76:44 CpuInfo.scala 77:10]
  always @(posedge clock) begin
    masterReg_Cmd <= io_ocp_M_Cmd; // @[CpuInfo.scala 26:22]
    masterReg_Addr <= io_ocp_M_Addr; // @[CpuInfo.scala 26:22]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  masterReg_Cmd = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  masterReg_Addr = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Leds(
  input         clock,
  input         reset,
  input  [2:0]  io_ocp_M_Cmd,
  input  [31:0] io_ocp_M_Data,
  output [1:0]  io_ocp_S_Resp,
  output [31:0] io_ocp_S_Data,
  output [8:0]  io_pins_led
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] ledReg; // @[Leds.scala 34:19]
  reg [1:0] respReg; // @[Leds.scala 37:20]
  reg [8:0] REG; // @[Leds.scala 56:21]
  assign io_ocp_S_Resp = respReg; // @[Leds.scala 52:17]
  assign io_ocp_S_Data = {{23'd0}, ledReg}; // @[Leds.scala 53:17]
  assign io_pins_led = REG; // @[Leds.scala 56:15]
  always @(posedge clock) begin
    if (reset) begin // @[Leds.scala 34:19]
      ledReg <= 9'h0; // @[Leds.scala 34:19]
    end else if (io_ocp_M_Cmd == 3'h1) begin // @[Leds.scala 41:36]
      ledReg <= io_ocp_M_Data[8:0]; // @[Leds.scala 43:12]
    end
    if (reset) begin // @[Leds.scala 37:20]
      respReg <= 2'h0; // @[Leds.scala 37:20]
    end else if (io_ocp_M_Cmd == 3'h2) begin // @[Leds.scala 47:36]
      respReg <= 2'h1; // @[Leds.scala 48:13]
    end else if (io_ocp_M_Cmd == 3'h1) begin // @[Leds.scala 41:36]
      respReg <= 2'h1; // @[Leds.scala 42:13]
    end else begin
      respReg <= 2'h0; // @[Leds.scala 38:11]
    end
    REG <= ledReg; // @[Leds.scala 56:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ledReg = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  respReg = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  REG = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Keys(
  input         clock,
  input         reset,
  input  [2:0]  io_ocp_M_Cmd,
  output [1:0]  io_ocp_S_Resp,
  output [31:0] io_ocp_S_Data,
  input  [3:0]  io_pins_key,
  output        io_interrupts_0,
  output        io_interrupts_1,
  output        io_interrupts_2,
  output        io_interrupts_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] keySyncReg; // @[Keys.scala 35:23]
  reg [3:0] keyReg; // @[Keys.scala 36:19]
  reg [1:0] respReg; // @[Keys.scala 39:20]
  assign io_ocp_S_Resp = respReg; // @[Keys.scala 48:17]
  assign io_ocp_S_Data = {{28'd0}, keyReg}; // @[Keys.scala 49:17]
  assign io_interrupts_0 = keyReg[0] & ~keySyncReg[0]; // @[Keys.scala 57:50]
  assign io_interrupts_1 = keyReg[1] & ~keySyncReg[1]; // @[Keys.scala 57:50]
  assign io_interrupts_2 = keyReg[2] & ~keySyncReg[2]; // @[Keys.scala 57:50]
  assign io_interrupts_3 = keyReg[3] & ~keySyncReg[3]; // @[Keys.scala 57:50]
  always @(posedge clock) begin
    keySyncReg <= io_pins_key; // @[Keys.scala 52:14]
    keyReg <= keySyncReg; // @[Keys.scala 53:10]
    if (reset) begin // @[Keys.scala 39:20]
      respReg <= 2'h0; // @[Keys.scala 39:20]
    end else if (io_ocp_M_Cmd == 3'h2) begin // @[Keys.scala 43:36]
      respReg <= 2'h1; // @[Keys.scala 44:13]
    end else begin
      respReg <= 2'h0; // @[Keys.scala 40:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  keySyncReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  keyReg = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  respReg = _RAND_2[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Timer(
  input         clock,
  input         reset,
  input  [2:0]  io_ocp_M_Cmd,
  input  [31:0] io_ocp_M_Addr,
  input  [31:0] io_ocp_M_Data,
  output [1:0]  io_ocp_S_Resp,
  output [31:0] io_ocp_S_Data,
  output        io_interrupts_0,
  output        io_interrupts_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] masterReg_Cmd; // @[Timer.scala 32:22]
  reg [31:0] masterReg_Addr; // @[Timer.scala 32:22]
  reg [31:0] masterReg_Data; // @[Timer.scala 32:22]
  reg [63:0] cycleReg; // @[Timer.scala 35:25]
  reg [63:0] cycleIntrReg; // @[Timer.scala 36:25]
  reg [6:0] usecSubReg; // @[Timer.scala 40:24]
  reg [63:0] usecReg; // @[Timer.scala 41:24]
  reg [63:0] usecIntrReg; // @[Timer.scala 42:24]
  reg [31:0] cycleHiReg; // @[Timer.scala 45:24]
  reg [31:0] usecHiReg; // @[Timer.scala 46:24]
  reg [31:0] cycleLoReg; // @[Timer.scala 49:24]
  reg [31:0] usecLoReg; // @[Timer.scala 50:24]
  wire  _T_2 = masterReg_Addr[3:2] == 2'h1; // @[Timer.scala 64:31]
  wire [31:0] _GEN_0 = masterReg_Addr[3:2] == 2'h1 ? cycleReg[31:0] : 32'h0; // @[Timer.scala 64:48 Timer.scala 65:12 Timer.scala 56:8]
  wire  _T_6 = masterReg_Addr[3:2] == 2'h0; // @[Timer.scala 68:31]
  wire [31:0] _GEN_2 = masterReg_Addr[3:2] == 2'h0 ? cycleHiReg : _GEN_0; // @[Timer.scala 68:48 Timer.scala 69:12]
  wire  _T_8 = masterReg_Addr[3:2] == 2'h3; // @[Timer.scala 74:31]
  wire [31:0] _GEN_3 = masterReg_Addr[3:2] == 2'h3 ? usecReg[31:0] : _GEN_2; // @[Timer.scala 74:48 Timer.scala 75:12]
  wire  _T_12 = masterReg_Addr[3:2] == 2'h2; // @[Timer.scala 78:31]
  wire [31:0] _GEN_5 = masterReg_Addr[3:2] == 2'h2 ? usecHiReg : _GEN_3; // @[Timer.scala 78:48 Timer.scala 79:12]
  wire [1:0] _GEN_6 = masterReg_Cmd == 3'h2 ? 2'h1 : 2'h0; // @[Timer.scala 59:37 Timer.scala 60:10 Timer.scala 55:8]
  wire [63:0] _T_18 = {masterReg_Data,cycleLoReg}; // @[Timer.scala 93:38]
  wire [63:0] _T_23 = {masterReg_Data,usecLoReg}; // @[Timer.scala 102:37]
  wire [63:0] _T_25 = cycleReg + 64'h1; // @[Timer.scala 115:24]
  wire [6:0] _T_30 = usecSubReg + 7'h1; // @[Timer.scala 121:28]
  wire [6:0] _T_32 = 7'h50 - 7'h1; // @[Timer.scala 122:34]
  wire [63:0] _T_35 = usecReg + 64'h1; // @[Timer.scala 124:24]
  wire  _T_38 = _T_35 == usecIntrReg; // @[Timer.scala 126:29]
  assign io_ocp_S_Resp = masterReg_Cmd == 3'h1 ? 2'h1 : _GEN_6; // @[Timer.scala 84:37 Timer.scala 85:10]
  assign io_ocp_S_Data = masterReg_Cmd == 3'h2 ? _GEN_5 : 32'h0; // @[Timer.scala 59:37 Timer.scala 56:8]
  assign io_interrupts_0 = _T_25 == cycleIntrReg; // @[Timer.scala 117:28]
  assign io_interrupts_1 = usecSubReg == _T_32 & _T_38; // @[Timer.scala 122:45 Timer.scala 112:20]
  always @(posedge clock) begin
    masterReg_Cmd <= io_ocp_M_Cmd; // @[Timer.scala 32:22]
    masterReg_Addr <= io_ocp_M_Addr; // @[Timer.scala 32:22]
    masterReg_Data <= io_ocp_M_Data; // @[Timer.scala 32:22]
    if (reset) begin // @[Timer.scala 35:25]
      cycleReg <= 64'h0; // @[Timer.scala 35:25]
    end else begin
      cycleReg <= _T_25; // @[Timer.scala 115:12]
    end
    if (reset) begin // @[Timer.scala 36:25]
      cycleIntrReg <= 64'h0; // @[Timer.scala 36:25]
    end else if (masterReg_Cmd == 3'h1) begin // @[Timer.scala 84:37]
      if (_T_6) begin // @[Timer.scala 92:48]
        cycleIntrReg <= _T_18; // @[Timer.scala 93:20]
      end
    end
    if (reset) begin // @[Timer.scala 40:24]
      usecSubReg <= 7'h0; // @[Timer.scala 40:24]
    end else if (usecSubReg == _T_32) begin // @[Timer.scala 122:45]
      usecSubReg <= 7'h0; // @[Timer.scala 123:16]
    end else begin
      usecSubReg <= _T_30; // @[Timer.scala 121:14]
    end
    if (reset) begin // @[Timer.scala 41:24]
      usecReg <= 64'h0; // @[Timer.scala 41:24]
    end else if (usecSubReg == _T_32) begin // @[Timer.scala 122:45]
      usecReg <= _T_35; // @[Timer.scala 124:13]
    end
    if (reset) begin // @[Timer.scala 42:24]
      usecIntrReg <= 64'h0; // @[Timer.scala 42:24]
    end else if (masterReg_Cmd == 3'h1) begin // @[Timer.scala 84:37]
      if (_T_12) begin // @[Timer.scala 101:48]
        usecIntrReg <= _T_23; // @[Timer.scala 102:19]
      end
    end
    if (masterReg_Cmd == 3'h2) begin // @[Timer.scala 59:37]
      if (masterReg_Addr[3:2] == 2'h1) begin // @[Timer.scala 64:48]
        cycleHiReg <= cycleReg[63:32]; // @[Timer.scala 66:18]
      end
    end
    if (masterReg_Cmd == 3'h2) begin // @[Timer.scala 59:37]
      if (masterReg_Addr[3:2] == 2'h3) begin // @[Timer.scala 74:48]
        usecHiReg <= usecReg[63:32]; // @[Timer.scala 76:17]
      end
    end
    if (masterReg_Cmd == 3'h1) begin // @[Timer.scala 84:37]
      if (_T_2) begin // @[Timer.scala 89:48]
        cycleLoReg <= masterReg_Data; // @[Timer.scala 90:18]
      end
    end
    if (masterReg_Cmd == 3'h1) begin // @[Timer.scala 84:37]
      if (_T_8) begin // @[Timer.scala 98:48]
        usecLoReg <= masterReg_Data; // @[Timer.scala 99:17]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  masterReg_Cmd = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  masterReg_Addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  masterReg_Data = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  cycleReg = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  cycleIntrReg = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  usecSubReg = _RAND_5[6:0];
  _RAND_6 = {2{`RANDOM}};
  usecReg = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  usecIntrReg = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  cycleHiReg = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  usecHiReg = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  cycleLoReg = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  usecLoReg = _RAND_11[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Deadline(
  input         clock,
  input         reset,
  input  [2:0]  io_ocp_M_Cmd,
  input  [31:0] io_ocp_M_Data,
  output [1:0]  io_ocp_S_Resp,
  output [31:0] io_ocp_S_Data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] downCountReg; // @[Deadline.scala 65:25]
  wire  downDone = downCountReg == 32'h0; // @[Deadline.scala 68:31]
  wire  _T_2 = ~downDone; // @[Deadline.scala 70:9]
  wire [31:0] _T_4 = downCountReg - 32'h1; // @[Deadline.scala 71:34]
  wire  _T_5 = io_ocp_M_Cmd == 3'h1; // @[Deadline.scala 73:22]
  reg  stallReg; // @[Deadline.scala 78:21]
  reg [1:0] respReg; // @[Deadline.scala 83:20]
  wire  _T_6 = io_ocp_M_Cmd == 3'h2; // @[Deadline.scala 86:22]
  wire  _GEN_3 = _T_6 & _T_2 | stallReg; // @[Deadline.scala 90:52 Deadline.scala 91:14 Deadline.scala 78:21]
  assign io_ocp_S_Resp = respReg; // @[Deadline.scala 101:17]
  assign io_ocp_S_Data = downCountReg; // @[Deadline.scala 100:17]
  always @(posedge clock) begin
    if (reset) begin // @[Deadline.scala 65:25]
      downCountReg <= 32'h0; // @[Deadline.scala 65:25]
    end else if (io_ocp_M_Cmd == 3'h1) begin // @[Deadline.scala 73:37]
      downCountReg <= io_ocp_M_Data; // @[Deadline.scala 74:18]
    end else if (~downDone) begin // @[Deadline.scala 70:20]
      downCountReg <= _T_4; // @[Deadline.scala 71:18]
    end
    if (reset) begin // @[Deadline.scala 78:21]
      stallReg <= 1'h0; // @[Deadline.scala 78:21]
    end else if (stallReg & downDone) begin // @[Deadline.scala 95:31]
      stallReg <= 1'h0; // @[Deadline.scala 97:14]
    end else begin
      stallReg <= _GEN_3;
    end
    if (reset) begin // @[Deadline.scala 83:20]
      respReg <= 2'h0; // @[Deadline.scala 83:20]
    end else if (stallReg & downDone) begin // @[Deadline.scala 95:31]
      respReg <= 2'h1; // @[Deadline.scala 96:13]
    end else if (io_ocp_M_Cmd == 3'h2 & downDone | _T_5) begin // @[Deadline.scala 86:80]
      respReg <= 2'h1; // @[Deadline.scala 87:13]
    end else begin
      respReg <= 2'h0; // @[Deadline.scala 84:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  downCountReg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  stallReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  respReg = _RAND_2[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Spm(
  input         clock,
  input  [2:0]  io_M_Cmd,
  input  [10:0] io_M_Addr,
  input  [31:0] io_M_Data,
  input  [3:0]  io_M_ByteEn,
  output [1:0]  io_S_Resp,
  output [31:0] io_S_Data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  MemBlock_clock; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_io_rdData; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_io_wrData; // @[MemBlock.scala 15:11]
  wire  MemBlock_1_clock; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_1_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_1_io_rdData; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_1_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_1_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_1_io_wrData; // @[MemBlock.scala 15:11]
  wire  MemBlock_2_clock; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_2_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_2_io_rdData; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_2_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_2_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_2_io_wrData; // @[MemBlock.scala 15:11]
  wire  MemBlock_3_clock; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_3_io_rdAddr; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_3_io_rdData; // @[MemBlock.scala 15:11]
  wire [8:0] MemBlock_3_io_wrAddr; // @[MemBlock.scala 15:11]
  wire  MemBlock_3_io_wrEna; // @[MemBlock.scala 15:11]
  wire [7:0] MemBlock_3_io_wrData; // @[MemBlock.scala 15:11]
  reg [2:0] cmdReg; // @[Spm.scala 32:19]
  wire [3:0] _T_5 = io_M_Cmd == 3'h1 ? io_M_ByteEn : 4'h0; // @[Spm.scala 45:20]
  wire [23:0] _T_23 = {MemBlock_2_io_rdData,MemBlock_1_io_rdData,MemBlock_io_rdData}; // @[Spm.scala 52:79]
  MemBlock_9 MemBlock ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_clock),
    .io_rdAddr(MemBlock_io_rdAddr),
    .io_rdData(MemBlock_io_rdData),
    .io_wrAddr(MemBlock_io_wrAddr),
    .io_wrEna(MemBlock_io_wrEna),
    .io_wrData(MemBlock_io_wrData)
  );
  MemBlock_9 MemBlock_1 ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_1_clock),
    .io_rdAddr(MemBlock_1_io_rdAddr),
    .io_rdData(MemBlock_1_io_rdData),
    .io_wrAddr(MemBlock_1_io_wrAddr),
    .io_wrEna(MemBlock_1_io_wrEna),
    .io_wrData(MemBlock_1_io_wrData)
  );
  MemBlock_9 MemBlock_2 ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_2_clock),
    .io_rdAddr(MemBlock_2_io_rdAddr),
    .io_rdData(MemBlock_2_io_rdData),
    .io_wrAddr(MemBlock_2_io_wrAddr),
    .io_wrEna(MemBlock_2_io_wrEna),
    .io_wrData(MemBlock_2_io_wrData)
  );
  MemBlock_9 MemBlock_3 ( // @[MemBlock.scala 15:11]
    .clock(MemBlock_3_clock),
    .io_rdAddr(MemBlock_3_io_rdAddr),
    .io_rdData(MemBlock_3_io_rdData),
    .io_wrAddr(MemBlock_3_io_wrAddr),
    .io_wrEna(MemBlock_3_io_wrEna),
    .io_wrData(MemBlock_3_io_wrData)
  );
  assign io_S_Resp = cmdReg == 3'h1 | cmdReg == 3'h2 ? 2'h1 : 2'h0; // @[Spm.scala 33:19]
  assign io_S_Data = {MemBlock_3_io_rdData,_T_23}; // @[Spm.scala 52:79]
  assign MemBlock_clock = clock;
  assign MemBlock_io_rdAddr = io_M_Addr[10:2]; // @[Spm.scala 52:37]
  assign MemBlock_io_wrAddr = io_M_Addr[10:2]; // @[Spm.scala 47:37]
  assign MemBlock_io_wrEna = _T_5[0]; // @[Spm.scala 47:23]
  assign MemBlock_io_wrData = io_M_Data[7:0]; // @[Spm.scala 48:27]
  assign MemBlock_1_clock = clock;
  assign MemBlock_1_io_rdAddr = io_M_Addr[10:2]; // @[Spm.scala 52:37]
  assign MemBlock_1_io_wrAddr = io_M_Addr[10:2]; // @[Spm.scala 47:37]
  assign MemBlock_1_io_wrEna = _T_5[1]; // @[Spm.scala 47:23]
  assign MemBlock_1_io_wrData = io_M_Data[15:8]; // @[Spm.scala 48:27]
  assign MemBlock_2_clock = clock;
  assign MemBlock_2_io_rdAddr = io_M_Addr[10:2]; // @[Spm.scala 52:37]
  assign MemBlock_2_io_wrAddr = io_M_Addr[10:2]; // @[Spm.scala 47:37]
  assign MemBlock_2_io_wrEna = _T_5[2]; // @[Spm.scala 47:23]
  assign MemBlock_2_io_wrData = io_M_Data[23:16]; // @[Spm.scala 48:27]
  assign MemBlock_3_clock = clock;
  assign MemBlock_3_io_rdAddr = io_M_Addr[10:2]; // @[Spm.scala 52:37]
  assign MemBlock_3_io_wrAddr = io_M_Addr[10:2]; // @[Spm.scala 47:37]
  assign MemBlock_3_io_wrEna = _T_5[3]; // @[Spm.scala 47:23]
  assign MemBlock_3_io_wrData = io_M_Data[31:24]; // @[Spm.scala 48:27]
  always @(posedge clock) begin
    cmdReg <= io_M_Cmd; // @[Spm.scala 32:19]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cmdReg = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SRamCtrl(
  input         clock,
  input         reset,
  input  [2:0]  io_ocp_M_Cmd,
  input  [20:0] io_ocp_M_Addr,
  input  [31:0] io_ocp_M_Data,
  input         io_ocp_M_DataValid,
  input  [3:0]  io_ocp_M_DataByteEn,
  output [1:0]  io_ocp_S_Resp,
  output [31:0] io_ocp_S_Data,
  output [19:0] io_pins_ramOut_addr,
  output        io_pins_ramOut_doutEna,
  output [15:0] io_pins_ramOut_dout,
  output        io_pins_ramOut_noe,
  output        io_pins_ramOut_nwe,
  output        io_pins_ramOut_nlb,
  output        io_pins_ramOut_nub,
  input  [15:0] io_pins_ramIn_din
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] stateReg; // @[SRamCtrl.scala 80:21]
  reg [19:0] mAddrReg; // @[SRamCtrl.scala 83:21]
  reg [15:0] rdBufferReg_0; // @[SRamCtrl.scala 84:24]
  reg [15:0] rdBufferReg_1; // @[SRamCtrl.scala 84:24]
  reg [15:0] rdBufferReg_2; // @[SRamCtrl.scala 84:24]
  reg [15:0] rdBufferReg_3; // @[SRamCtrl.scala 84:24]
  reg [15:0] rdBufferReg_4; // @[SRamCtrl.scala 84:24]
  reg [15:0] rdBufferReg_5; // @[SRamCtrl.scala 84:24]
  reg [15:0] rdBufferReg_6; // @[SRamCtrl.scala 84:24]
  reg [15:0] rdBufferReg_7; // @[SRamCtrl.scala 84:24]
  reg [1:0] wrBufferReg_0_byteEna; // @[SRamCtrl.scala 85:24]
  reg [15:0] wrBufferReg_0_data; // @[SRamCtrl.scala 85:24]
  reg [1:0] wrBufferReg_1_byteEna; // @[SRamCtrl.scala 85:24]
  reg [15:0] wrBufferReg_1_data; // @[SRamCtrl.scala 85:24]
  reg [1:0] wrBufferReg_2_byteEna; // @[SRamCtrl.scala 85:24]
  reg [15:0] wrBufferReg_2_data; // @[SRamCtrl.scala 85:24]
  reg [1:0] wrBufferReg_3_byteEna; // @[SRamCtrl.scala 85:24]
  reg [15:0] wrBufferReg_3_data; // @[SRamCtrl.scala 85:24]
  reg [1:0] wrBufferReg_4_byteEna; // @[SRamCtrl.scala 85:24]
  reg [15:0] wrBufferReg_4_data; // @[SRamCtrl.scala 85:24]
  reg [1:0] wrBufferReg_5_byteEna; // @[SRamCtrl.scala 85:24]
  reg [15:0] wrBufferReg_5_data; // @[SRamCtrl.scala 85:24]
  reg [1:0] wrBufferReg_6_byteEna; // @[SRamCtrl.scala 85:24]
  reg [15:0] wrBufferReg_6_data; // @[SRamCtrl.scala 85:24]
  reg [1:0] wrBufferReg_7_byteEna; // @[SRamCtrl.scala 85:24]
  reg [15:0] wrBufferReg_7_data; // @[SRamCtrl.scala 85:24]
  reg [2:0] transCountReg; // @[SRamCtrl.scala 86:26]
  reg [1:0] wordCountReg; // @[SRamCtrl.scala 87:25]
  reg  waitCountReg; // @[SRamCtrl.scala 88:25]
  reg [19:0] addrReg; // @[SRamCtrl.scala 90:20]
  reg  doutEnaReg; // @[SRamCtrl.scala 91:23]
  reg [31:0] doutReg; // @[SRamCtrl.scala 92:20]
  reg  noeReg; // @[SRamCtrl.scala 94:19]
  reg  nweReg; // @[SRamCtrl.scala 95:19]
  reg  nlbReg; // @[SRamCtrl.scala 96:19]
  reg  nubReg; // @[SRamCtrl.scala 97:19]
  wire [2:0] _T_9 = {wordCountReg,1'h0}; // @[SRamCtrl.scala 104:45]
  wire [2:0] _T_10 = {wordCountReg,1'h1}; // @[SRamCtrl.scala 104:45]
  wire [15:0] _GEN_1 = 3'h1 == _T_10 ? rdBufferReg_1 : rdBufferReg_0; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_2 = 3'h2 == _T_10 ? rdBufferReg_2 : _GEN_1; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_3 = 3'h3 == _T_10 ? rdBufferReg_3 : _GEN_2; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_4 = 3'h4 == _T_10 ? rdBufferReg_4 : _GEN_3; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_5 = 3'h5 == _T_10 ? rdBufferReg_5 : _GEN_4; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_6 = 3'h6 == _T_10 ? rdBufferReg_6 : _GEN_5; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_7 = 3'h7 == _T_10 ? rdBufferReg_7 : _GEN_6; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_9 = 3'h1 == _T_9 ? rdBufferReg_1 : rdBufferReg_0; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_10 = 3'h2 == _T_9 ? rdBufferReg_2 : _GEN_9; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_11 = 3'h3 == _T_9 ? rdBufferReg_3 : _GEN_10; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_12 = 3'h4 == _T_9 ? rdBufferReg_4 : _GEN_11; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_13 = 3'h5 == _T_9 ? rdBufferReg_5 : _GEN_12; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_14 = 3'h6 == _T_9 ? rdBufferReg_6 : _GEN_13; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [15:0] _GEN_15 = 3'h7 == _T_9 ? rdBufferReg_7 : _GEN_14; // @[SRamCtrl.scala 105:47 SRamCtrl.scala 105:47]
  wire [2:0] _GEN_16 = io_ocp_M_Cmd == 3'h2 ? 3'h1 : stateReg; // @[SRamCtrl.scala 127:40 SRamCtrl.scala 128:18 SRamCtrl.scala 80:21]
  wire [1:0] _GEN_17 = io_ocp_M_Cmd == 3'h1 ? 2'h1 : wordCountReg; // @[SRamCtrl.scala 130:40 SRamCtrl.scala 131:22 SRamCtrl.scala 87:25]
  wire [2:0] _GEN_18 = io_ocp_M_Cmd == 3'h1 ? 3'h4 : _GEN_16; // @[SRamCtrl.scala 130:40 SRamCtrl.scala 132:18]
  wire [19:0] _GEN_19 = io_ocp_M_Cmd != 3'h0 ? io_ocp_M_Addr[20:1] : mAddrReg; // @[SRamCtrl.scala 124:40 SRamCtrl.scala 125:16 SRamCtrl.scala 83:21]
  wire [2:0] _GEN_20 = io_ocp_M_Cmd != 3'h0 ? _GEN_18 : stateReg; // @[SRamCtrl.scala 124:40 SRamCtrl.scala 80:21]
  wire [1:0] _GEN_21 = io_ocp_M_Cmd != 3'h0 ? _GEN_17 : wordCountReg; // @[SRamCtrl.scala 124:40 SRamCtrl.scala 87:25]
  wire [1:0] _GEN_22 = stateReg == 3'h0 ? io_ocp_M_DataByteEn[1:0] : wrBufferReg_0_byteEna; // @[SRamCtrl.scala 119:29 SRamCtrl.scala 121:30 SRamCtrl.scala 85:24]
  wire [15:0] _GEN_23 = stateReg == 3'h0 ? io_ocp_M_Data[15:0] : wrBufferReg_0_data; // @[SRamCtrl.scala 119:29 SRamCtrl.scala 122:27 SRamCtrl.scala 85:24]
  wire [1:0] _GEN_24 = stateReg == 3'h0 ? io_ocp_M_DataByteEn[3:2] : wrBufferReg_1_byteEna; // @[SRamCtrl.scala 119:29 SRamCtrl.scala 121:30 SRamCtrl.scala 85:24]
  wire [15:0] _GEN_25 = stateReg == 3'h0 ? io_ocp_M_Data[31:16] : wrBufferReg_1_data; // @[SRamCtrl.scala 119:29 SRamCtrl.scala 122:27 SRamCtrl.scala 85:24]
  wire [19:0] _GEN_26 = stateReg == 3'h0 ? _GEN_19 : mAddrReg; // @[SRamCtrl.scala 119:29 SRamCtrl.scala 83:21]
  wire [2:0] _GEN_27 = stateReg == 3'h0 ? _GEN_20 : stateReg; // @[SRamCtrl.scala 119:29 SRamCtrl.scala 80:21]
  wire [1:0] _GEN_28 = stateReg == 3'h0 ? _GEN_21 : wordCountReg; // @[SRamCtrl.scala 119:29 SRamCtrl.scala 87:25]
  wire  _GEN_29 = stateReg == 3'h1 ? 1'h0 : 1'h1; // @[SRamCtrl.scala 136:31 SRamCtrl.scala 137:12 SRamCtrl.scala 112:10]
  wire [2:0] _GEN_31 = stateReg == 3'h1 ? 3'h2 : _GEN_27; // @[SRamCtrl.scala 136:31 SRamCtrl.scala 153:16]
  wire [19:0] _T_24 = mAddrReg + 20'h1; // @[SRamCtrl.scala 161:25]
  wire [2:0] _T_28 = transCountReg + 3'h1; // @[SRamCtrl.scala 165:36]
  wire  _T_29 = transCountReg == 3'h7; // @[SRamCtrl.scala 167:24]
  wire [2:0] _GEN_32 = transCountReg == 3'h7 ? 3'h3 : 3'h1; // @[SRamCtrl.scala 167:48 SRamCtrl.scala 168:16 SRamCtrl.scala 166:14]
  wire [2:0] _GEN_33 = transCountReg == 3'h7 ? 3'h0 : _T_28; // @[SRamCtrl.scala 167:48 SRamCtrl.scala 169:21 SRamCtrl.scala 165:19]
  wire  _GEN_34 = stateReg == 3'h2 ? 1'h0 : _GEN_29; // @[SRamCtrl.scala 156:32 SRamCtrl.scala 157:12]
  wire [19:0] _GEN_36 = stateReg == 3'h2 ? _T_24 : mAddrReg; // @[SRamCtrl.scala 156:32 SRamCtrl.scala 161:13 SRamCtrl.scala 108:11]
  wire [19:0] _GEN_37 = stateReg == 3'h2 ? _T_24 : _GEN_26; // @[SRamCtrl.scala 156:32 SRamCtrl.scala 162:14]
  wire [2:0] _GEN_46 = stateReg == 3'h2 ? _GEN_33 : transCountReg; // @[SRamCtrl.scala 156:32 SRamCtrl.scala 86:26]
  wire [2:0] _GEN_47 = stateReg == 3'h2 ? _GEN_32 : _GEN_31; // @[SRamCtrl.scala 156:32]
  wire [1:0] _T_32 = wordCountReg + 2'h1; // @[SRamCtrl.scala 174:34]
  wire  _T_33 = wordCountReg == 2'h3; // @[SRamCtrl.scala 175:23]
  wire [2:0] _GEN_48 = wordCountReg == 2'h3 ? 3'h0 : _GEN_47; // @[SRamCtrl.scala 175:47 SRamCtrl.scala 176:16]
  wire [1:0] _GEN_49 = wordCountReg == 2'h3 ? 2'h0 : _T_32; // @[SRamCtrl.scala 175:47 SRamCtrl.scala 177:20 SRamCtrl.scala 174:18]
  wire [1:0] _GEN_50 = stateReg == 3'h3 ? 2'h1 : 2'h0; // @[SRamCtrl.scala 172:31 SRamCtrl.scala 173:19 SRamCtrl.scala 100:17]
  wire [1:0] _GEN_51 = stateReg == 3'h3 ? _GEN_49 : _GEN_28; // @[SRamCtrl.scala 172:31]
  wire [2:0] _GEN_52 = stateReg == 3'h3 ? _GEN_48 : _GEN_47; // @[SRamCtrl.scala 172:31]
  wire  _T_34 = stateReg == 3'h4; // @[SRamCtrl.scala 180:17]
  wire [2:0] _GEN_85 = _T_33 ? 3'h5 : _GEN_52; // @[SRamCtrl.scala 191:49 SRamCtrl.scala 192:18]
  wire [2:0] _GEN_89 = io_ocp_M_DataValid ? _GEN_85 : 3'h4; // @[SRamCtrl.scala 189:41 SRamCtrl.scala 197:16]
  wire  _GEN_90 = io_ocp_M_DataValid & _T_33; // @[SRamCtrl.scala 189:41 SRamCtrl.scala 117:16]
  wire  _GEN_92 = _T_33 ? 1'h0 : 1'h1; // @[SRamCtrl.scala 199:47 SRamCtrl.scala 201:14 SRamCtrl.scala 113:10]
  wire  _GEN_93 = _T_33 ? ~wrBufferReg_0_byteEna[1] : _GEN_34; // @[SRamCtrl.scala 199:47 SRamCtrl.scala 202:14]
  wire  _GEN_94 = _T_33 ? ~wrBufferReg_0_byteEna[0] : _GEN_34; // @[SRamCtrl.scala 199:47 SRamCtrl.scala 203:14]
  wire [2:0] _GEN_114 = stateReg == 3'h4 ? _GEN_89 : _GEN_52; // @[SRamCtrl.scala 180:32]
  wire  _GEN_115 = stateReg == 3'h4 & _GEN_90; // @[SRamCtrl.scala 180:32 SRamCtrl.scala 117:16]
  wire  _GEN_117 = stateReg == 3'h4 ? _GEN_92 : 1'h1; // @[SRamCtrl.scala 180:32 SRamCtrl.scala 113:10]
  wire  _GEN_118 = stateReg == 3'h4 ? _GEN_93 : _GEN_34; // @[SRamCtrl.scala 180:32]
  wire  _GEN_119 = stateReg == 3'h4 ? _GEN_94 : _GEN_34; // @[SRamCtrl.scala 180:32]
  wire [1:0] _GEN_122 = 3'h1 == transCountReg ? wrBufferReg_1_byteEna : wrBufferReg_0_byteEna; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [15:0] _GEN_123 = 3'h1 == transCountReg ? wrBufferReg_1_data : wrBufferReg_0_data; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [1:0] _GEN_124 = 3'h2 == transCountReg ? wrBufferReg_2_byteEna : _GEN_122; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [15:0] _GEN_125 = 3'h2 == transCountReg ? wrBufferReg_2_data : _GEN_123; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [1:0] _GEN_126 = 3'h3 == transCountReg ? wrBufferReg_3_byteEna : _GEN_124; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [15:0] _GEN_127 = 3'h3 == transCountReg ? wrBufferReg_3_data : _GEN_125; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [1:0] _GEN_128 = 3'h4 == transCountReg ? wrBufferReg_4_byteEna : _GEN_126; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [15:0] _GEN_129 = 3'h4 == transCountReg ? wrBufferReg_4_data : _GEN_127; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [1:0] _GEN_130 = 3'h5 == transCountReg ? wrBufferReg_5_byteEna : _GEN_128; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [15:0] _GEN_131 = 3'h5 == transCountReg ? wrBufferReg_5_data : _GEN_129; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [1:0] _GEN_132 = 3'h6 == transCountReg ? wrBufferReg_6_byteEna : _GEN_130; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [15:0] _GEN_133 = 3'h6 == transCountReg ? wrBufferReg_6_data : _GEN_131; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [1:0] _GEN_134 = 3'h7 == transCountReg ? wrBufferReg_7_byteEna : _GEN_132; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire [15:0] _GEN_135 = 3'h7 == transCountReg ? wrBufferReg_7_data : _GEN_133; // @[SRamCtrl.scala 209:13 SRamCtrl.scala 209:13]
  wire  _GEN_136 = waitCountReg < 1'h1 & waitCountReg + 1'h1; // @[SRamCtrl.scala 211:47 SRamCtrl.scala 212:20 SRamCtrl.scala 217:20]
  wire  _GEN_137 = waitCountReg < 1'h1 ? ~_GEN_134[1] : 1'h1; // @[SRamCtrl.scala 211:47 SRamCtrl.scala 213:14 SRamCtrl.scala 218:14]
  wire  _GEN_138 = waitCountReg < 1'h1 ? ~_GEN_134[0] : 1'h1; // @[SRamCtrl.scala 211:47 SRamCtrl.scala 214:14 SRamCtrl.scala 219:14]
  wire [2:0] _GEN_139 = waitCountReg < 1'h1 ? 3'h5 : 3'h6; // @[SRamCtrl.scala 211:47 SRamCtrl.scala 215:16 SRamCtrl.scala 220:16]
  wire  _GEN_141 = stateReg == 3'h5 ? 1'h0 : _GEN_117; // @[SRamCtrl.scala 206:32 SRamCtrl.scala 208:12]
  wire [15:0] _GEN_142 = stateReg == 3'h5 ? _GEN_135 : wrBufferReg_0_data; // @[SRamCtrl.scala 206:32 SRamCtrl.scala 209:13]
  wire  _GEN_143 = stateReg == 3'h5 | _T_34; // @[SRamCtrl.scala 206:32 SRamCtrl.scala 210:16]
  wire  _GEN_144 = stateReg == 3'h5 ? _GEN_136 : _GEN_115; // @[SRamCtrl.scala 206:32]
  wire  _GEN_145 = stateReg == 3'h5 ? _GEN_137 : _GEN_118; // @[SRamCtrl.scala 206:32]
  wire  _GEN_146 = stateReg == 3'h5 ? _GEN_138 : _GEN_119; // @[SRamCtrl.scala 206:32]
  wire [2:0] _GEN_147 = stateReg == 3'h5 ? _GEN_139 : _GEN_114; // @[SRamCtrl.scala 206:32]
  wire [1:0] _GEN_150 = 3'h1 == _T_28 ? wrBufferReg_1_byteEna : wrBufferReg_0_byteEna; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [15:0] _GEN_151 = 3'h1 == _T_28 ? wrBufferReg_1_data : wrBufferReg_0_data; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [1:0] _GEN_152 = 3'h2 == _T_28 ? wrBufferReg_2_byteEna : _GEN_150; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [15:0] _GEN_153 = 3'h2 == _T_28 ? wrBufferReg_2_data : _GEN_151; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [1:0] _GEN_154 = 3'h3 == _T_28 ? wrBufferReg_3_byteEna : _GEN_152; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [15:0] _GEN_155 = 3'h3 == _T_28 ? wrBufferReg_3_data : _GEN_153; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [1:0] _GEN_156 = 3'h4 == _T_28 ? wrBufferReg_4_byteEna : _GEN_154; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [15:0] _GEN_157 = 3'h4 == _T_28 ? wrBufferReg_4_data : _GEN_155; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [1:0] _GEN_158 = 3'h5 == _T_28 ? wrBufferReg_5_byteEna : _GEN_156; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [15:0] _GEN_159 = 3'h5 == _T_28 ? wrBufferReg_5_data : _GEN_157; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [1:0] _GEN_160 = 3'h6 == _T_28 ? wrBufferReg_6_byteEna : _GEN_158; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [15:0] _GEN_161 = 3'h6 == _T_28 ? wrBufferReg_6_data : _GEN_159; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [1:0] _GEN_162 = 3'h7 == _T_28 ? wrBufferReg_7_byteEna : _GEN_160; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [15:0] _GEN_163 = 3'h7 == _T_28 ? wrBufferReg_7_data : _GEN_161; // @[SRamCtrl.scala 227:60 SRamCtrl.scala 227:60]
  wire [15:0] _GEN_200 = transCountReg < 3'h7 ? _GEN_163 : _GEN_142; // @[SRamCtrl.scala 224:46 SRamCtrl.scala 229:15]
  wire  _GEN_201 = transCountReg < 3'h7 | _GEN_143; // @[SRamCtrl.scala 224:46 SRamCtrl.scala 230:18]
  wire  _GEN_205 = transCountReg < 3'h7 | _GEN_144; // @[SRamCtrl.scala 224:46 SRamCtrl.scala 234:20]
  wire [2:0] _GEN_206 = transCountReg < 3'h7 ? 3'h5 : _GEN_147; // @[SRamCtrl.scala 224:46 SRamCtrl.scala 235:16]
  wire [15:0] _GEN_214 = stateReg == 3'h6 ? _GEN_200 : _GEN_142; // @[SRamCtrl.scala 223:33]
  assign io_ocp_S_Resp = stateReg == 3'h7 ? 2'h1 : _GEN_50; // @[SRamCtrl.scala 243:32 SRamCtrl.scala 244:19]
  assign io_ocp_S_Data = {_GEN_7,_GEN_15}; // @[SRamCtrl.scala 105:47]
  assign io_pins_ramOut_addr = addrReg; // @[SRamCtrl.scala 248:23]
  assign io_pins_ramOut_doutEna = doutEnaReg; // @[SRamCtrl.scala 249:26]
  assign io_pins_ramOut_dout = doutReg[15:0]; // @[SRamCtrl.scala 250:23]
  assign io_pins_ramOut_noe = noeReg; // @[SRamCtrl.scala 252:22]
  assign io_pins_ramOut_nwe = nweReg; // @[SRamCtrl.scala 253:22]
  assign io_pins_ramOut_nlb = nlbReg; // @[SRamCtrl.scala 254:22]
  assign io_pins_ramOut_nub = nubReg; // @[SRamCtrl.scala 255:22]
  always @(posedge clock) begin
    if (reset) begin // @[SRamCtrl.scala 80:21]
      stateReg <= 3'h0; // @[SRamCtrl.scala 80:21]
    end else if (stateReg == 3'h7) begin // @[SRamCtrl.scala 243:32]
      stateReg <= 3'h0; // @[SRamCtrl.scala 245:14]
    end else if (stateReg == 3'h6) begin // @[SRamCtrl.scala 223:33]
      if (_T_29) begin // @[SRamCtrl.scala 237:48]
        stateReg <= 3'h7; // @[SRamCtrl.scala 238:16]
      end else begin
        stateReg <= _GEN_206;
      end
    end else if (stateReg == 3'h5) begin // @[SRamCtrl.scala 206:32]
      stateReg <= _GEN_139;
    end else begin
      stateReg <= _GEN_114;
    end
    if (stateReg == 3'h6) begin // @[SRamCtrl.scala 223:33]
      if (transCountReg < 3'h7) begin // @[SRamCtrl.scala 224:46]
        mAddrReg <= _T_24; // @[SRamCtrl.scala 232:16]
      end else begin
        mAddrReg <= _GEN_37;
      end
    end else begin
      mAddrReg <= _GEN_37;
    end
    if (stateReg == 3'h2) begin // @[SRamCtrl.scala 156:32]
      rdBufferReg_0 <= rdBufferReg_1; // @[SRamCtrl.scala 163:55]
    end
    if (stateReg == 3'h2) begin // @[SRamCtrl.scala 156:32]
      rdBufferReg_1 <= rdBufferReg_2; // @[SRamCtrl.scala 163:55]
    end
    if (stateReg == 3'h2) begin // @[SRamCtrl.scala 156:32]
      rdBufferReg_2 <= rdBufferReg_3; // @[SRamCtrl.scala 163:55]
    end
    if (stateReg == 3'h2) begin // @[SRamCtrl.scala 156:32]
      rdBufferReg_3 <= rdBufferReg_4; // @[SRamCtrl.scala 163:55]
    end
    if (stateReg == 3'h2) begin // @[SRamCtrl.scala 156:32]
      rdBufferReg_4 <= rdBufferReg_5; // @[SRamCtrl.scala 163:55]
    end
    if (stateReg == 3'h2) begin // @[SRamCtrl.scala 156:32]
      rdBufferReg_5 <= rdBufferReg_6; // @[SRamCtrl.scala 163:55]
    end
    if (stateReg == 3'h2) begin // @[SRamCtrl.scala 156:32]
      rdBufferReg_6 <= rdBufferReg_7; // @[SRamCtrl.scala 163:55]
    end
    if (stateReg == 3'h2) begin // @[SRamCtrl.scala 156:32]
      rdBufferReg_7 <= io_pins_ramIn_din; // @[SRamCtrl.scala 164:32]
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h0 == _T_10) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_0_byteEna <= io_ocp_M_DataByteEn[3:2]; // @[SRamCtrl.scala 182:52]
      end else if (3'h0 == _T_9) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_0_byteEna <= io_ocp_M_DataByteEn[1:0]; // @[SRamCtrl.scala 182:52]
      end else begin
        wrBufferReg_0_byteEna <= _GEN_22;
      end
    end else begin
      wrBufferReg_0_byteEna <= _GEN_22;
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h0 == _T_10) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_0_data <= io_ocp_M_Data[31:16]; // @[SRamCtrl.scala 184:49]
      end else if (3'h0 == _T_9) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_0_data <= io_ocp_M_Data[15:0]; // @[SRamCtrl.scala 184:49]
      end else begin
        wrBufferReg_0_data <= _GEN_23;
      end
    end else begin
      wrBufferReg_0_data <= _GEN_23;
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h1 == _T_10) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_1_byteEna <= io_ocp_M_DataByteEn[3:2]; // @[SRamCtrl.scala 182:52]
      end else if (3'h1 == _T_9) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_1_byteEna <= io_ocp_M_DataByteEn[1:0]; // @[SRamCtrl.scala 182:52]
      end else begin
        wrBufferReg_1_byteEna <= _GEN_24;
      end
    end else begin
      wrBufferReg_1_byteEna <= _GEN_24;
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h1 == _T_10) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_1_data <= io_ocp_M_Data[31:16]; // @[SRamCtrl.scala 184:49]
      end else if (3'h1 == _T_9) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_1_data <= io_ocp_M_Data[15:0]; // @[SRamCtrl.scala 184:49]
      end else begin
        wrBufferReg_1_data <= _GEN_25;
      end
    end else begin
      wrBufferReg_1_data <= _GEN_25;
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h2 == _T_10) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_2_byteEna <= io_ocp_M_DataByteEn[3:2]; // @[SRamCtrl.scala 182:52]
      end else if (3'h2 == _T_9) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_2_byteEna <= io_ocp_M_DataByteEn[1:0]; // @[SRamCtrl.scala 182:52]
      end
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h2 == _T_10) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_2_data <= io_ocp_M_Data[31:16]; // @[SRamCtrl.scala 184:49]
      end else if (3'h2 == _T_9) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_2_data <= io_ocp_M_Data[15:0]; // @[SRamCtrl.scala 184:49]
      end
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h3 == _T_10) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_3_byteEna <= io_ocp_M_DataByteEn[3:2]; // @[SRamCtrl.scala 182:52]
      end else if (3'h3 == _T_9) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_3_byteEna <= io_ocp_M_DataByteEn[1:0]; // @[SRamCtrl.scala 182:52]
      end
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h3 == _T_10) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_3_data <= io_ocp_M_Data[31:16]; // @[SRamCtrl.scala 184:49]
      end else if (3'h3 == _T_9) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_3_data <= io_ocp_M_Data[15:0]; // @[SRamCtrl.scala 184:49]
      end
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h4 == _T_10) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_4_byteEna <= io_ocp_M_DataByteEn[3:2]; // @[SRamCtrl.scala 182:52]
      end else if (3'h4 == _T_9) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_4_byteEna <= io_ocp_M_DataByteEn[1:0]; // @[SRamCtrl.scala 182:52]
      end
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h4 == _T_10) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_4_data <= io_ocp_M_Data[31:16]; // @[SRamCtrl.scala 184:49]
      end else if (3'h4 == _T_9) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_4_data <= io_ocp_M_Data[15:0]; // @[SRamCtrl.scala 184:49]
      end
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h5 == _T_10) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_5_byteEna <= io_ocp_M_DataByteEn[3:2]; // @[SRamCtrl.scala 182:52]
      end else if (3'h5 == _T_9) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_5_byteEna <= io_ocp_M_DataByteEn[1:0]; // @[SRamCtrl.scala 182:52]
      end
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h5 == _T_10) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_5_data <= io_ocp_M_Data[31:16]; // @[SRamCtrl.scala 184:49]
      end else if (3'h5 == _T_9) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_5_data <= io_ocp_M_Data[15:0]; // @[SRamCtrl.scala 184:49]
      end
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h6 == _T_10) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_6_byteEna <= io_ocp_M_DataByteEn[3:2]; // @[SRamCtrl.scala 182:52]
      end else if (3'h6 == _T_9) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_6_byteEna <= io_ocp_M_DataByteEn[1:0]; // @[SRamCtrl.scala 182:52]
      end
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h6 == _T_10) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_6_data <= io_ocp_M_Data[31:16]; // @[SRamCtrl.scala 184:49]
      end else if (3'h6 == _T_9) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_6_data <= io_ocp_M_Data[15:0]; // @[SRamCtrl.scala 184:49]
      end
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h7 == _T_10) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_7_byteEna <= io_ocp_M_DataByteEn[3:2]; // @[SRamCtrl.scala 182:52]
      end else if (3'h7 == _T_9) begin // @[SRamCtrl.scala 182:52]
        wrBufferReg_7_byteEna <= io_ocp_M_DataByteEn[1:0]; // @[SRamCtrl.scala 182:52]
      end
    end
    if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (3'h7 == _T_10) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_7_data <= io_ocp_M_Data[31:16]; // @[SRamCtrl.scala 184:49]
      end else if (3'h7 == _T_9) begin // @[SRamCtrl.scala 184:49]
        wrBufferReg_7_data <= io_ocp_M_Data[15:0]; // @[SRamCtrl.scala 184:49]
      end
    end
    if (reset) begin // @[SRamCtrl.scala 86:26]
      transCountReg <= 3'h0; // @[SRamCtrl.scala 86:26]
    end else if (stateReg == 3'h6) begin // @[SRamCtrl.scala 223:33]
      if (_T_29) begin // @[SRamCtrl.scala 237:48]
        transCountReg <= 3'h0; // @[SRamCtrl.scala 239:21]
      end else if (transCountReg < 3'h7) begin // @[SRamCtrl.scala 224:46]
        transCountReg <= _T_28; // @[SRamCtrl.scala 233:21]
      end else begin
        transCountReg <= _GEN_46;
      end
    end else begin
      transCountReg <= _GEN_46;
    end
    if (reset) begin // @[SRamCtrl.scala 87:25]
      wordCountReg <= 2'h0; // @[SRamCtrl.scala 87:25]
    end else if (stateReg == 3'h4) begin // @[SRamCtrl.scala 180:32]
      if (io_ocp_M_DataValid) begin // @[SRamCtrl.scala 189:41]
        wordCountReg <= _GEN_49;
      end else begin
        wordCountReg <= _GEN_51;
      end
    end else begin
      wordCountReg <= _GEN_51;
    end
    if (reset) begin // @[SRamCtrl.scala 88:25]
      waitCountReg <= 1'h0; // @[SRamCtrl.scala 88:25]
    end else if (stateReg == 3'h6) begin // @[SRamCtrl.scala 223:33]
      if (_T_29) begin // @[SRamCtrl.scala 237:48]
        waitCountReg <= 1'h0; // @[SRamCtrl.scala 240:20]
      end else begin
        waitCountReg <= _GEN_205;
      end
    end else if (stateReg == 3'h5) begin // @[SRamCtrl.scala 206:32]
      waitCountReg <= _GEN_136;
    end else begin
      waitCountReg <= _GEN_115;
    end
    if (stateReg == 3'h6) begin // @[SRamCtrl.scala 223:33]
      if (transCountReg < 3'h7) begin // @[SRamCtrl.scala 224:46]
        addrReg <= _T_24; // @[SRamCtrl.scala 231:15]
      end else begin
        addrReg <= _GEN_36;
      end
    end else begin
      addrReg <= _GEN_36;
    end
    if (stateReg == 3'h6) begin // @[SRamCtrl.scala 223:33]
      doutEnaReg <= _GEN_201;
    end else begin
      doutEnaReg <= _GEN_143;
    end
    doutReg <= {{16'd0}, _GEN_214}; // @[SRamCtrl.scala 223:33]
    if (stateReg == 3'h2) begin // @[SRamCtrl.scala 156:32]
      noeReg <= 1'h0; // @[SRamCtrl.scala 157:12]
    end else if (stateReg == 3'h1) begin // @[SRamCtrl.scala 136:31]
      noeReg <= 1'h0; // @[SRamCtrl.scala 137:12]
    end else begin
      noeReg <= 1'h1; // @[SRamCtrl.scala 112:10]
    end
    if (stateReg == 3'h6) begin // @[SRamCtrl.scala 223:33]
      if (transCountReg < 3'h7) begin // @[SRamCtrl.scala 224:46]
        nweReg <= 1'h0; // @[SRamCtrl.scala 226:14]
      end else begin
        nweReg <= _GEN_141;
      end
    end else begin
      nweReg <= _GEN_141;
    end
    if (stateReg == 3'h6) begin // @[SRamCtrl.scala 223:33]
      if (transCountReg < 3'h7) begin // @[SRamCtrl.scala 224:46]
        nlbReg <= ~_GEN_162[0]; // @[SRamCtrl.scala 228:14]
      end else begin
        nlbReg <= _GEN_146;
      end
    end else begin
      nlbReg <= _GEN_146;
    end
    if (stateReg == 3'h6) begin // @[SRamCtrl.scala 223:33]
      if (transCountReg < 3'h7) begin // @[SRamCtrl.scala 224:46]
        nubReg <= ~_GEN_162[1]; // @[SRamCtrl.scala 227:14]
      end else begin
        nubReg <= _GEN_145;
      end
    end else begin
      nubReg <= _GEN_145;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  mAddrReg = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  rdBufferReg_0 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  rdBufferReg_1 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  rdBufferReg_2 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  rdBufferReg_3 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  rdBufferReg_4 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  rdBufferReg_5 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  rdBufferReg_6 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  rdBufferReg_7 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  wrBufferReg_0_byteEna = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  wrBufferReg_0_data = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  wrBufferReg_1_byteEna = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  wrBufferReg_1_data = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  wrBufferReg_2_byteEna = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  wrBufferReg_2_data = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  wrBufferReg_3_byteEna = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  wrBufferReg_3_data = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  wrBufferReg_4_byteEna = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  wrBufferReg_4_data = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  wrBufferReg_5_byteEna = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  wrBufferReg_5_data = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  wrBufferReg_6_byteEna = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  wrBufferReg_6_data = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  wrBufferReg_7_byteEna = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  wrBufferReg_7_data = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  transCountReg = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  wordCountReg = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  waitCountReg = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  addrReg = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  doutEnaReg = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  doutReg = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  noeReg = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  nweReg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  nlbReg = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  nubReg = _RAND_35[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Patmos(
  input         clock,
  input         reset,
  output [8:0]  io_Leds_led,
  output        io_UartCmp_tx,
  output [19:0] io_SRamCtrl_ramOut_addr,
  output        io_SRamCtrl_ramOut_doutEna,
  output [15:0] io_SRamCtrl_ramOut_dout,
  output        io_SRamCtrl_ramOut_nce,
  output        io_SRamCtrl_ramOut_noe,
  output        io_SRamCtrl_ramOut_nwe,
  output        io_SRamCtrl_ramOut_nlb,
  output        io_SRamCtrl_ramOut_nub,
  input  [3:0]  io_Keys_key,
  input         io_UartCmp_rx,
  input  [15:0] io_SRamCtrl_ramIn_din
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  cores_0_clock; // @[Patmos.scala 213:48]
  wire  cores_0_reset; // @[Patmos.scala 213:48]
  wire  cores_0_io_interrupts_0; // @[Patmos.scala 213:48]
  wire  cores_0_io_interrupts_1; // @[Patmos.scala 213:48]
  wire  cores_0_io_interrupts_2; // @[Patmos.scala 213:48]
  wire  cores_0_io_interrupts_3; // @[Patmos.scala 213:48]
  wire  cores_0_io_interrupts_4; // @[Patmos.scala 213:48]
  wire  cores_0_io_interrupts_5; // @[Patmos.scala 213:48]
  wire [2:0] cores_0_io_memPort_M_Cmd; // @[Patmos.scala 213:48]
  wire [20:0] cores_0_io_memPort_M_Addr; // @[Patmos.scala 213:48]
  wire [31:0] cores_0_io_memPort_M_Data; // @[Patmos.scala 213:48]
  wire  cores_0_io_memPort_M_DataValid; // @[Patmos.scala 213:48]
  wire [3:0] cores_0_io_memPort_M_DataByteEn; // @[Patmos.scala 213:48]
  wire [1:0] cores_0_io_memPort_S_Resp; // @[Patmos.scala 213:48]
  wire [31:0] cores_0_io_memPort_S_Data; // @[Patmos.scala 213:48]
  wire [2:0] cores_0_io_memInOut_M_Cmd; // @[Patmos.scala 213:48]
  wire [31:0] cores_0_io_memInOut_M_Addr; // @[Patmos.scala 213:48]
  wire [31:0] cores_0_io_memInOut_M_Data; // @[Patmos.scala 213:48]
  wire [3:0] cores_0_io_memInOut_M_ByteEn; // @[Patmos.scala 213:48]
  wire [1:0] cores_0_io_memInOut_S_Resp; // @[Patmos.scala 213:48]
  wire [31:0] cores_0_io_memInOut_S_Data; // @[Patmos.scala 213:48]
  wire [2:0] cores_0_io_excInOut_M_Cmd; // @[Patmos.scala 213:48]
  wire [31:0] cores_0_io_excInOut_M_Addr; // @[Patmos.scala 213:48]
  wire [31:0] cores_0_io_excInOut_M_Data; // @[Patmos.scala 213:48]
  wire [1:0] cores_0_io_excInOut_S_Resp; // @[Patmos.scala 213:48]
  wire [31:0] cores_0_io_excInOut_S_Data; // @[Patmos.scala 213:48]
  wire  HardlockOCPWrapper_clock; // @[Patmos.scala 248:63]
  wire  HardlockOCPWrapper_reset; // @[Patmos.scala 248:63]
  wire [2:0] HardlockOCPWrapper_io_cores_0_M_Cmd; // @[Patmos.scala 248:63]
  wire [1:0] HardlockOCPWrapper_io_cores_0_S_Resp; // @[Patmos.scala 248:63]
  wire  UartCmp_clock; // @[Patmos.scala 257:62]
  wire  UartCmp_reset; // @[Patmos.scala 257:62]
  wire [2:0] UartCmp_io_cores_0_M_Cmd; // @[Patmos.scala 257:62]
  wire [31:0] UartCmp_io_cores_0_M_Addr; // @[Patmos.scala 257:62]
  wire [31:0] UartCmp_io_cores_0_M_Data; // @[Patmos.scala 257:62]
  wire [1:0] UartCmp_io_cores_0_S_Resp; // @[Patmos.scala 257:62]
  wire [31:0] UartCmp_io_cores_0_S_Data; // @[Patmos.scala 257:62]
  wire  UartCmp_io_pins_tx; // @[Patmos.scala 257:62]
  wire  UartCmp_io_pins_rx; // @[Patmos.scala 257:62]
  wire  CpuInfo_clock; // @[Patmos.scala 282:25]
  wire [2:0] CpuInfo_io_ocp_M_Cmd; // @[Patmos.scala 282:25]
  wire [31:0] CpuInfo_io_ocp_M_Addr; // @[Patmos.scala 282:25]
  wire [1:0] CpuInfo_io_ocp_S_Resp; // @[Patmos.scala 282:25]
  wire [31:0] CpuInfo_io_ocp_S_Data; // @[Patmos.scala 282:25]
  wire  Leds_clock; // @[Leds.scala 22:11]
  wire  Leds_reset; // @[Leds.scala 22:11]
  wire [2:0] Leds_io_ocp_M_Cmd; // @[Leds.scala 22:11]
  wire [31:0] Leds_io_ocp_M_Data; // @[Leds.scala 22:11]
  wire [1:0] Leds_io_ocp_S_Resp; // @[Leds.scala 22:11]
  wire [31:0] Leds_io_ocp_S_Data; // @[Leds.scala 22:11]
  wire [8:0] Leds_io_pins_led; // @[Leds.scala 22:11]
  wire  Keys_clock; // @[Keys.scala 22:11]
  wire  Keys_reset; // @[Keys.scala 22:11]
  wire [2:0] Keys_io_ocp_M_Cmd; // @[Keys.scala 22:11]
  wire [1:0] Keys_io_ocp_S_Resp; // @[Keys.scala 22:11]
  wire [31:0] Keys_io_ocp_S_Data; // @[Keys.scala 22:11]
  wire [3:0] Keys_io_pins_key; // @[Keys.scala 22:11]
  wire  Keys_io_interrupts_0; // @[Keys.scala 22:11]
  wire  Keys_io_interrupts_1; // @[Keys.scala 22:11]
  wire  Keys_io_interrupts_2; // @[Keys.scala 22:11]
  wire  Keys_io_interrupts_3; // @[Keys.scala 22:11]
  wire  Timer_clock; // @[Timer.scala 22:11]
  wire  Timer_reset; // @[Timer.scala 22:11]
  wire [2:0] Timer_io_ocp_M_Cmd; // @[Timer.scala 22:11]
  wire [31:0] Timer_io_ocp_M_Addr; // @[Timer.scala 22:11]
  wire [31:0] Timer_io_ocp_M_Data; // @[Timer.scala 22:11]
  wire [1:0] Timer_io_ocp_S_Resp; // @[Timer.scala 22:11]
  wire [31:0] Timer_io_ocp_S_Data; // @[Timer.scala 22:11]
  wire  Timer_io_interrupts_0; // @[Timer.scala 22:11]
  wire  Timer_io_interrupts_1; // @[Timer.scala 22:11]
  wire  Deadline_clock; // @[Deadline.scala 53:61]
  wire  Deadline_reset; // @[Deadline.scala 53:61]
  wire [2:0] Deadline_io_ocp_M_Cmd; // @[Deadline.scala 53:61]
  wire [31:0] Deadline_io_ocp_M_Data; // @[Deadline.scala 53:61]
  wire [1:0] Deadline_io_ocp_S_Resp; // @[Deadline.scala 53:61]
  wire [31:0] Deadline_io_ocp_S_Data; // @[Deadline.scala 53:61]
  wire  Spm_clock; // @[Patmos.scala 335:21]
  wire [2:0] Spm_io_M_Cmd; // @[Patmos.scala 335:21]
  wire [10:0] Spm_io_M_Addr; // @[Patmos.scala 335:21]
  wire [31:0] Spm_io_M_Data; // @[Patmos.scala 335:21]
  wire [3:0] Spm_io_M_ByteEn; // @[Patmos.scala 335:21]
  wire [1:0] Spm_io_S_Resp; // @[Patmos.scala 335:21]
  wire [31:0] Spm_io_S_Data; // @[Patmos.scala 335:21]
  wire  ramCtrl_clock; // @[SRamCtrl.scala 34:11]
  wire  ramCtrl_reset; // @[SRamCtrl.scala 34:11]
  wire [2:0] ramCtrl_io_ocp_M_Cmd; // @[SRamCtrl.scala 34:11]
  wire [20:0] ramCtrl_io_ocp_M_Addr; // @[SRamCtrl.scala 34:11]
  wire [31:0] ramCtrl_io_ocp_M_Data; // @[SRamCtrl.scala 34:11]
  wire  ramCtrl_io_ocp_M_DataValid; // @[SRamCtrl.scala 34:11]
  wire [3:0] ramCtrl_io_ocp_M_DataByteEn; // @[SRamCtrl.scala 34:11]
  wire [1:0] ramCtrl_io_ocp_S_Resp; // @[SRamCtrl.scala 34:11]
  wire [31:0] ramCtrl_io_ocp_S_Data; // @[SRamCtrl.scala 34:11]
  wire [19:0] ramCtrl_io_pins_ramOut_addr; // @[SRamCtrl.scala 34:11]
  wire  ramCtrl_io_pins_ramOut_doutEna; // @[SRamCtrl.scala 34:11]
  wire [15:0] ramCtrl_io_pins_ramOut_dout; // @[SRamCtrl.scala 34:11]
  wire  ramCtrl_io_pins_ramOut_noe; // @[SRamCtrl.scala 34:11]
  wire  ramCtrl_io_pins_ramOut_nwe; // @[SRamCtrl.scala 34:11]
  wire  ramCtrl_io_pins_ramOut_nlb; // @[SRamCtrl.scala 34:11]
  wire  ramCtrl_io_pins_ramOut_nub; // @[SRamCtrl.scala 34:11]
  wire [15:0] ramCtrl_io_pins_ramIn_din; // @[SRamCtrl.scala 34:11]
  wire  _T_41 = cores_0_io_memInOut_M_Addr[31:16] == 16'h1; // @[Patmos.scala 385:85]
  wire [2:0] _GEN_36 = _T_41 ? cores_0_io_memInOut_M_Cmd : 3'h0; // @[Patmos.scala 390:17 Patmos.scala 391:19 Patmos.scala 389:17]
  reg [1:0] REG; // @[Patmos.scala 340:29]
  wire  _T_3 = cores_0_io_memInOut_M_Addr[31:16] == 16'hf009; // @[Patmos.scala 385:85]
  reg  REG_1; // @[Patmos.scala 394:27]
  wire  _T_5 = cores_0_io_memInOut_M_Cmd != 3'h0; // @[Patmos.scala 395:39]
  wire [31:0] _GEN_3 = REG_1 ? Leds_io_ocp_S_Data : 32'h0; // @[Patmos.scala 398:20 Patmos.scala 399:37 Patmos.scala 379:33]
  wire  _T_7 = cores_0_io_memInOut_M_Addr[31:16] == 16'hf00a; // @[Patmos.scala 385:85]
  reg  REG_2; // @[Patmos.scala 394:27]
  wire [31:0] _GEN_7 = REG_2 ? Keys_io_ocp_S_Data : _GEN_3; // @[Patmos.scala 398:20 Patmos.scala 399:37]
  wire  _T_11 = cores_0_io_memInOut_M_Addr[31:16] == 16'hf002; // @[Patmos.scala 385:85]
  reg  REG_3; // @[Patmos.scala 394:27]
  wire [31:0] _GEN_11 = REG_3 ? Timer_io_ocp_S_Data : _GEN_7; // @[Patmos.scala 398:20 Patmos.scala 399:37]
  wire  _T_15 = cores_0_io_memInOut_M_Addr[31:16] == 16'hf003; // @[Patmos.scala 385:85]
  reg  REG_4; // @[Patmos.scala 394:27]
  wire [31:0] _GEN_15 = REG_4 ? Deadline_io_ocp_S_Data : _GEN_11; // @[Patmos.scala 398:20 Patmos.scala 399:37]
  wire  _T_19 = cores_0_io_memInOut_M_Addr[31:16] == 16'hf000; // @[Patmos.scala 385:85]
  reg  REG_5; // @[Patmos.scala 394:27]
  wire [31:0] _GEN_19 = REG_5 ? CpuInfo_io_ocp_S_Data : _GEN_15; // @[Patmos.scala 398:20 Patmos.scala 399:37]
  wire  _T_23 = cores_0_io_memInOut_M_Addr[31:16] == 16'hf001; // @[Patmos.scala 385:85]
  reg  REG_6; // @[Patmos.scala 394:27]
  wire [31:0] _GEN_23 = REG_6 ? cores_0_io_excInOut_S_Data : _GEN_19; // @[Patmos.scala 398:20 Patmos.scala 399:37]
  wire  _T_27 = cores_0_io_memInOut_M_Addr[31:16] == 16'he801; // @[Patmos.scala 385:85]
  reg  REG_7; // @[Patmos.scala 394:27]
  wire [31:0] _GEN_27 = REG_7 ? 32'h0 : _GEN_23; // @[Patmos.scala 398:20 Patmos.scala 399:37]
  wire  _T_31 = cores_0_io_memInOut_M_Addr[31:16] == 16'hf008; // @[Patmos.scala 385:85]
  reg  REG_8; // @[Patmos.scala 394:27]
  wire [31:0] _GEN_31 = REG_8 ? UartCmp_io_cores_0_S_Data : _GEN_27; // @[Patmos.scala 398:20 Patmos.scala 399:37]
  wire  _T_37 = ~cores_0_io_memInOut_M_Addr[16]; // @[Patmos.scala 386:32]
  wire  _T_38 = cores_0_io_memInOut_M_Addr[31:28] == 4'h0 & _T_37; // @[Patmos.scala 385:100]
  reg  REG_9; // @[Patmos.scala 394:27]
  wire [31:0] _GEN_35 = REG_9 ? Spm_io_S_Data : _GEN_31; // @[Patmos.scala 398:20 Patmos.scala 399:37]
  wire  _GEN_37 = _T_41 | (_T_38 | (_T_31 | (_T_27 | (_T_23 | (_T_19 | (_T_15 | (_T_11 | (_T_7 | _T_3)))))))); // @[Patmos.scala 390:17 Patmos.scala 392:18]
  reg  REG_10; // @[Patmos.scala 394:27]
  reg [1:0] REG_11; // @[Patmos.scala 418:25]
  wire [1:0] _T_47 = Leds_io_ocp_S_Resp; // @[Patmos.scala 424:122]
  wire [1:0] _T_48 = _T_47 | Keys_io_ocp_S_Resp; // @[Patmos.scala 424:122]
  wire [1:0] _T_49 = _T_48 | Timer_io_ocp_S_Resp; // @[Patmos.scala 424:122]
  wire [1:0] _T_50 = _T_49 | Deadline_io_ocp_S_Resp; // @[Patmos.scala 424:122]
  wire [1:0] _T_51 = _T_50 | CpuInfo_io_ocp_S_Resp; // @[Patmos.scala 424:122]
  wire [1:0] _T_52 = _T_51 | cores_0_io_excInOut_S_Resp; // @[Patmos.scala 424:122]
  wire [1:0] _T_53 = _T_52 | HardlockOCPWrapper_io_cores_0_S_Resp; // @[Patmos.scala 424:122]
  wire [1:0] _T_54 = _T_53 | UartCmp_io_cores_0_S_Resp; // @[Patmos.scala 424:122]
  wire [1:0] _T_55 = _T_54 | Spm_io_S_Resp; // @[Patmos.scala 424:122]
  wire [1:0] _T_56 = _T_55 | REG; // @[Patmos.scala 424:122]
  PatmosCore cores_0 ( // @[Patmos.scala 213:48]
    .clock(cores_0_clock),
    .reset(cores_0_reset),
    .io_interrupts_0(cores_0_io_interrupts_0),
    .io_interrupts_1(cores_0_io_interrupts_1),
    .io_interrupts_2(cores_0_io_interrupts_2),
    .io_interrupts_3(cores_0_io_interrupts_3),
    .io_interrupts_4(cores_0_io_interrupts_4),
    .io_interrupts_5(cores_0_io_interrupts_5),
    .io_memPort_M_Cmd(cores_0_io_memPort_M_Cmd),
    .io_memPort_M_Addr(cores_0_io_memPort_M_Addr),
    .io_memPort_M_Data(cores_0_io_memPort_M_Data),
    .io_memPort_M_DataValid(cores_0_io_memPort_M_DataValid),
    .io_memPort_M_DataByteEn(cores_0_io_memPort_M_DataByteEn),
    .io_memPort_S_Resp(cores_0_io_memPort_S_Resp),
    .io_memPort_S_Data(cores_0_io_memPort_S_Data),
    .io_memInOut_M_Cmd(cores_0_io_memInOut_M_Cmd),
    .io_memInOut_M_Addr(cores_0_io_memInOut_M_Addr),
    .io_memInOut_M_Data(cores_0_io_memInOut_M_Data),
    .io_memInOut_M_ByteEn(cores_0_io_memInOut_M_ByteEn),
    .io_memInOut_S_Resp(cores_0_io_memInOut_S_Resp),
    .io_memInOut_S_Data(cores_0_io_memInOut_S_Data),
    .io_excInOut_M_Cmd(cores_0_io_excInOut_M_Cmd),
    .io_excInOut_M_Addr(cores_0_io_excInOut_M_Addr),
    .io_excInOut_M_Data(cores_0_io_excInOut_M_Data),
    .io_excInOut_S_Resp(cores_0_io_excInOut_S_Resp),
    .io_excInOut_S_Data(cores_0_io_excInOut_S_Data)
  );
  HardlockOCPWrapper HardlockOCPWrapper ( // @[Patmos.scala 248:63]
    .clock(HardlockOCPWrapper_clock),
    .reset(HardlockOCPWrapper_reset),
    .io_cores_0_M_Cmd(HardlockOCPWrapper_io_cores_0_M_Cmd),
    .io_cores_0_S_Resp(HardlockOCPWrapper_io_cores_0_S_Resp)
  );
  UartCmp UartCmp ( // @[Patmos.scala 257:62]
    .clock(UartCmp_clock),
    .reset(UartCmp_reset),
    .io_cores_0_M_Cmd(UartCmp_io_cores_0_M_Cmd),
    .io_cores_0_M_Addr(UartCmp_io_cores_0_M_Addr),
    .io_cores_0_M_Data(UartCmp_io_cores_0_M_Data),
    .io_cores_0_S_Resp(UartCmp_io_cores_0_S_Resp),
    .io_cores_0_S_Data(UartCmp_io_cores_0_S_Data),
    .io_pins_tx(UartCmp_io_pins_tx),
    .io_pins_rx(UartCmp_io_pins_rx)
  );
  CpuInfo CpuInfo ( // @[Patmos.scala 282:25]
    .clock(CpuInfo_clock),
    .io_ocp_M_Cmd(CpuInfo_io_ocp_M_Cmd),
    .io_ocp_M_Addr(CpuInfo_io_ocp_M_Addr),
    .io_ocp_S_Resp(CpuInfo_io_ocp_S_Resp),
    .io_ocp_S_Data(CpuInfo_io_ocp_S_Data)
  );
  Leds Leds ( // @[Leds.scala 22:11]
    .clock(Leds_clock),
    .reset(Leds_reset),
    .io_ocp_M_Cmd(Leds_io_ocp_M_Cmd),
    .io_ocp_M_Data(Leds_io_ocp_M_Data),
    .io_ocp_S_Resp(Leds_io_ocp_S_Resp),
    .io_ocp_S_Data(Leds_io_ocp_S_Data),
    .io_pins_led(Leds_io_pins_led)
  );
  Keys Keys ( // @[Keys.scala 22:11]
    .clock(Keys_clock),
    .reset(Keys_reset),
    .io_ocp_M_Cmd(Keys_io_ocp_M_Cmd),
    .io_ocp_S_Resp(Keys_io_ocp_S_Resp),
    .io_ocp_S_Data(Keys_io_ocp_S_Data),
    .io_pins_key(Keys_io_pins_key),
    .io_interrupts_0(Keys_io_interrupts_0),
    .io_interrupts_1(Keys_io_interrupts_1),
    .io_interrupts_2(Keys_io_interrupts_2),
    .io_interrupts_3(Keys_io_interrupts_3)
  );
  Timer Timer ( // @[Timer.scala 22:11]
    .clock(Timer_clock),
    .reset(Timer_reset),
    .io_ocp_M_Cmd(Timer_io_ocp_M_Cmd),
    .io_ocp_M_Addr(Timer_io_ocp_M_Addr),
    .io_ocp_M_Data(Timer_io_ocp_M_Data),
    .io_ocp_S_Resp(Timer_io_ocp_S_Resp),
    .io_ocp_S_Data(Timer_io_ocp_S_Data),
    .io_interrupts_0(Timer_io_interrupts_0),
    .io_interrupts_1(Timer_io_interrupts_1)
  );
  Deadline Deadline ( // @[Deadline.scala 53:61]
    .clock(Deadline_clock),
    .reset(Deadline_reset),
    .io_ocp_M_Cmd(Deadline_io_ocp_M_Cmd),
    .io_ocp_M_Data(Deadline_io_ocp_M_Data),
    .io_ocp_S_Resp(Deadline_io_ocp_S_Resp),
    .io_ocp_S_Data(Deadline_io_ocp_S_Data)
  );
  Spm Spm ( // @[Patmos.scala 335:21]
    .clock(Spm_clock),
    .io_M_Cmd(Spm_io_M_Cmd),
    .io_M_Addr(Spm_io_M_Addr),
    .io_M_Data(Spm_io_M_Data),
    .io_M_ByteEn(Spm_io_M_ByteEn),
    .io_S_Resp(Spm_io_S_Resp),
    .io_S_Data(Spm_io_S_Data)
  );
  SRamCtrl ramCtrl ( // @[SRamCtrl.scala 34:11]
    .clock(ramCtrl_clock),
    .reset(ramCtrl_reset),
    .io_ocp_M_Cmd(ramCtrl_io_ocp_M_Cmd),
    .io_ocp_M_Addr(ramCtrl_io_ocp_M_Addr),
    .io_ocp_M_Data(ramCtrl_io_ocp_M_Data),
    .io_ocp_M_DataValid(ramCtrl_io_ocp_M_DataValid),
    .io_ocp_M_DataByteEn(ramCtrl_io_ocp_M_DataByteEn),
    .io_ocp_S_Resp(ramCtrl_io_ocp_S_Resp),
    .io_ocp_S_Data(ramCtrl_io_ocp_S_Data),
    .io_pins_ramOut_addr(ramCtrl_io_pins_ramOut_addr),
    .io_pins_ramOut_doutEna(ramCtrl_io_pins_ramOut_doutEna),
    .io_pins_ramOut_dout(ramCtrl_io_pins_ramOut_dout),
    .io_pins_ramOut_noe(ramCtrl_io_pins_ramOut_noe),
    .io_pins_ramOut_nwe(ramCtrl_io_pins_ramOut_nwe),
    .io_pins_ramOut_nlb(ramCtrl_io_pins_ramOut_nlb),
    .io_pins_ramOut_nub(ramCtrl_io_pins_ramOut_nub),
    .io_pins_ramIn_din(ramCtrl_io_pins_ramIn_din)
  );
  assign io_Leds_led = Leds_io_pins_led; // @[Patmos.scala 461:36]
  assign io_UartCmp_tx = UartCmp_io_pins_tx; // @[Patmos.scala 461:36]
  assign io_SRamCtrl_ramOut_addr = ramCtrl_io_pins_ramOut_addr; // @[Patmos.scala 461:36]
  assign io_SRamCtrl_ramOut_doutEna = ramCtrl_io_pins_ramOut_doutEna; // @[Patmos.scala 461:36]
  assign io_SRamCtrl_ramOut_dout = ramCtrl_io_pins_ramOut_dout; // @[Patmos.scala 461:36]
  assign io_SRamCtrl_ramOut_nce = 1'h0; // @[Patmos.scala 461:36]
  assign io_SRamCtrl_ramOut_noe = ramCtrl_io_pins_ramOut_noe; // @[Patmos.scala 461:36]
  assign io_SRamCtrl_ramOut_nwe = ramCtrl_io_pins_ramOut_nwe; // @[Patmos.scala 461:36]
  assign io_SRamCtrl_ramOut_nlb = ramCtrl_io_pins_ramOut_nlb; // @[Patmos.scala 461:36]
  assign io_SRamCtrl_ramOut_nub = ramCtrl_io_pins_ramOut_nub; // @[Patmos.scala 461:36]
  assign cores_0_clock = clock;
  assign cores_0_reset = reset;
  assign cores_0_io_interrupts_0 = Timer_io_interrupts_0; // @[Patmos.scala 304:53]
  assign cores_0_io_interrupts_1 = Timer_io_interrupts_1; // @[Patmos.scala 304:53]
  assign cores_0_io_interrupts_2 = Keys_io_interrupts_0; // @[Patmos.scala 304:53]
  assign cores_0_io_interrupts_3 = Keys_io_interrupts_1; // @[Patmos.scala 304:53]
  assign cores_0_io_interrupts_4 = Keys_io_interrupts_2; // @[Patmos.scala 304:53]
  assign cores_0_io_interrupts_5 = Keys_io_interrupts_3; // @[Patmos.scala 304:53]
  assign cores_0_io_memPort_S_Resp = ramCtrl_io_ocp_S_Resp; // @[Patmos.scala 437:27]
  assign cores_0_io_memPort_S_Data = ramCtrl_io_ocp_S_Data; // @[Patmos.scala 437:27]
  assign cores_0_io_memInOut_S_Resp = REG_11 | _T_56; // @[Patmos.scala 424:47]
  assign cores_0_io_memInOut_S_Data = REG_10 ? 32'h0 : _GEN_35; // @[Patmos.scala 398:20 Patmos.scala 399:37]
  assign cores_0_io_excInOut_M_Cmd = _T_23 ? cores_0_io_memInOut_M_Cmd : 3'h0; // @[Patmos.scala 390:17 Patmos.scala 391:19 Patmos.scala 389:17]
  assign cores_0_io_excInOut_M_Addr = cores_0_io_memInOut_M_Addr; // @[Patmos.scala 388:13]
  assign cores_0_io_excInOut_M_Data = cores_0_io_memInOut_M_Data; // @[Patmos.scala 388:13]
  assign HardlockOCPWrapper_clock = clock;
  assign HardlockOCPWrapper_reset = reset;
  assign HardlockOCPWrapper_io_cores_0_M_Cmd = _T_27 ? cores_0_io_memInOut_M_Cmd : 3'h0; // @[Patmos.scala 390:17 Patmos.scala 391:19 Patmos.scala 389:17]
  assign UartCmp_clock = clock;
  assign UartCmp_reset = reset;
  assign UartCmp_io_cores_0_M_Cmd = _T_31 ? cores_0_io_memInOut_M_Cmd : 3'h0; // @[Patmos.scala 390:17 Patmos.scala 391:19 Patmos.scala 389:17]
  assign UartCmp_io_cores_0_M_Addr = cores_0_io_memInOut_M_Addr; // @[Patmos.scala 388:13]
  assign UartCmp_io_cores_0_M_Data = cores_0_io_memInOut_M_Data; // @[Patmos.scala 388:13]
  assign UartCmp_io_pins_rx = io_UartCmp_rx; // @[Patmos.scala 460:35]
  assign CpuInfo_clock = clock;
  assign CpuInfo_io_ocp_M_Cmd = _T_19 ? cores_0_io_memInOut_M_Cmd : 3'h0; // @[Patmos.scala 390:17 Patmos.scala 391:19 Patmos.scala 389:17]
  assign CpuInfo_io_ocp_M_Addr = cores_0_io_memInOut_M_Addr; // @[Patmos.scala 388:13]
  assign Leds_clock = clock;
  assign Leds_reset = reset;
  assign Leds_io_ocp_M_Cmd = _T_3 ? cores_0_io_memInOut_M_Cmd : 3'h0; // @[Patmos.scala 390:17 Patmos.scala 391:19 Patmos.scala 389:17]
  assign Leds_io_ocp_M_Data = cores_0_io_memInOut_M_Data; // @[Patmos.scala 388:13]
  assign Keys_clock = clock;
  assign Keys_reset = reset;
  assign Keys_io_ocp_M_Cmd = _T_7 ? cores_0_io_memInOut_M_Cmd : 3'h0; // @[Patmos.scala 390:17 Patmos.scala 391:19 Patmos.scala 389:17]
  assign Keys_io_pins_key = io_Keys_key; // @[Patmos.scala 460:35]
  assign Timer_clock = clock;
  assign Timer_reset = reset;
  assign Timer_io_ocp_M_Cmd = _T_11 ? cores_0_io_memInOut_M_Cmd : 3'h0; // @[Patmos.scala 390:17 Patmos.scala 391:19 Patmos.scala 389:17]
  assign Timer_io_ocp_M_Addr = cores_0_io_memInOut_M_Addr; // @[Patmos.scala 388:13]
  assign Timer_io_ocp_M_Data = cores_0_io_memInOut_M_Data; // @[Patmos.scala 388:13]
  assign Deadline_clock = clock;
  assign Deadline_reset = reset;
  assign Deadline_io_ocp_M_Cmd = _T_15 ? cores_0_io_memInOut_M_Cmd : 3'h0; // @[Patmos.scala 390:17 Patmos.scala 391:19 Patmos.scala 389:17]
  assign Deadline_io_ocp_M_Data = cores_0_io_memInOut_M_Data; // @[Patmos.scala 388:13]
  assign Spm_clock = clock;
  assign Spm_io_M_Cmd = _T_38 ? cores_0_io_memInOut_M_Cmd : 3'h0; // @[Patmos.scala 390:17 Patmos.scala 391:19 Patmos.scala 389:17]
  assign Spm_io_M_Addr = cores_0_io_memInOut_M_Addr[10:0]; // @[Patmos.scala 388:13]
  assign Spm_io_M_Data = cores_0_io_memInOut_M_Data; // @[Patmos.scala 388:13]
  assign Spm_io_M_ByteEn = cores_0_io_memInOut_M_ByteEn; // @[Patmos.scala 388:13]
  assign ramCtrl_clock = clock;
  assign ramCtrl_reset = reset;
  assign ramCtrl_io_ocp_M_Cmd = cores_0_io_memPort_M_Cmd; // @[Patmos.scala 436:22]
  assign ramCtrl_io_ocp_M_Addr = cores_0_io_memPort_M_Addr; // @[Patmos.scala 436:22]
  assign ramCtrl_io_ocp_M_Data = cores_0_io_memPort_M_Data; // @[Patmos.scala 436:22]
  assign ramCtrl_io_ocp_M_DataValid = cores_0_io_memPort_M_DataValid; // @[Patmos.scala 436:22]
  assign ramCtrl_io_ocp_M_DataByteEn = cores_0_io_memPort_M_DataByteEn; // @[Patmos.scala 436:22]
  assign ramCtrl_io_pins_ramIn_din = io_SRamCtrl_ramIn_din; // @[Patmos.scala 460:35]
  always @(posedge clock) begin
    if (_GEN_36 == 3'h0) begin // @[Patmos.scala 340:33]
      REG <= 2'h0;
    end else begin
      REG <= 2'h1;
    end
    if (reset) begin // @[Patmos.scala 394:27]
      REG_1 <= 1'h0; // @[Patmos.scala 394:27]
    end else if (cores_0_io_memInOut_M_Cmd != 3'h0) begin // @[Patmos.scala 395:56]
      REG_1 <= _T_3; // @[Patmos.scala 396:16]
    end
    if (reset) begin // @[Patmos.scala 394:27]
      REG_2 <= 1'h0; // @[Patmos.scala 394:27]
    end else if (cores_0_io_memInOut_M_Cmd != 3'h0) begin // @[Patmos.scala 395:56]
      REG_2 <= _T_7; // @[Patmos.scala 396:16]
    end
    if (reset) begin // @[Patmos.scala 394:27]
      REG_3 <= 1'h0; // @[Patmos.scala 394:27]
    end else if (cores_0_io_memInOut_M_Cmd != 3'h0) begin // @[Patmos.scala 395:56]
      REG_3 <= _T_11; // @[Patmos.scala 396:16]
    end
    if (reset) begin // @[Patmos.scala 394:27]
      REG_4 <= 1'h0; // @[Patmos.scala 394:27]
    end else if (cores_0_io_memInOut_M_Cmd != 3'h0) begin // @[Patmos.scala 395:56]
      REG_4 <= _T_15; // @[Patmos.scala 396:16]
    end
    if (reset) begin // @[Patmos.scala 394:27]
      REG_5 <= 1'h0; // @[Patmos.scala 394:27]
    end else if (cores_0_io_memInOut_M_Cmd != 3'h0) begin // @[Patmos.scala 395:56]
      REG_5 <= _T_19; // @[Patmos.scala 396:16]
    end
    if (reset) begin // @[Patmos.scala 394:27]
      REG_6 <= 1'h0; // @[Patmos.scala 394:27]
    end else if (cores_0_io_memInOut_M_Cmd != 3'h0) begin // @[Patmos.scala 395:56]
      REG_6 <= _T_23; // @[Patmos.scala 396:16]
    end
    if (reset) begin // @[Patmos.scala 394:27]
      REG_7 <= 1'h0; // @[Patmos.scala 394:27]
    end else if (cores_0_io_memInOut_M_Cmd != 3'h0) begin // @[Patmos.scala 395:56]
      REG_7 <= _T_27; // @[Patmos.scala 396:16]
    end
    if (reset) begin // @[Patmos.scala 394:27]
      REG_8 <= 1'h0; // @[Patmos.scala 394:27]
    end else if (cores_0_io_memInOut_M_Cmd != 3'h0) begin // @[Patmos.scala 395:56]
      REG_8 <= _T_31; // @[Patmos.scala 396:16]
    end
    if (reset) begin // @[Patmos.scala 394:27]
      REG_9 <= 1'h0; // @[Patmos.scala 394:27]
    end else if (cores_0_io_memInOut_M_Cmd != 3'h0) begin // @[Patmos.scala 395:56]
      REG_9 <= _T_38; // @[Patmos.scala 396:16]
    end
    if (reset) begin // @[Patmos.scala 394:27]
      REG_10 <= 1'h0; // @[Patmos.scala 394:27]
    end else if (cores_0_io_memInOut_M_Cmd != 3'h0) begin // @[Patmos.scala 395:56]
      REG_10 <= _T_41; // @[Patmos.scala 396:16]
    end
    if (reset) begin // @[Patmos.scala 418:25]
      REG_11 <= 2'h0; // @[Patmos.scala 418:25]
    end else if (_T_5 & ~_GEN_37) begin // @[Patmos.scala 419:67]
      REG_11 <= 2'h3; // @[Patmos.scala 420:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  REG_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  REG_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  REG_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG_11 = _RAND_11[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
